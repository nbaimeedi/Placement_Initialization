module gcd (clk,
    req_rdy,
    req_val,
    reset,
    resp_rdy,
    resp_val,
    req_msg,
    resp_msg);
 input clk;
 output req_rdy;
 input req_val;
 input reset;
 input resp_rdy;
 output resp_val;
 input [31:0] req_msg;
 output [15:0] resp_msg;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire \dpath.a_lt_b$in0[10] ;
 wire \dpath.a_lt_b$in0[11] ;
 wire \dpath.a_lt_b$in0[12] ;
 wire \dpath.a_lt_b$in0[13] ;
 wire \dpath.a_lt_b$in0[14] ;
 wire \dpath.a_lt_b$in0[15] ;
 wire \dpath.a_lt_b$in0[1] ;
 wire \dpath.a_lt_b$in0[2] ;
 wire \dpath.a_lt_b$in0[3] ;
 wire \dpath.a_lt_b$in0[4] ;
 wire \dpath.a_lt_b$in0[5] ;
 wire \dpath.a_lt_b$in0[6] ;
 wire \dpath.a_lt_b$in0[7] ;
 wire \dpath.a_lt_b$in0[8] ;
 wire \dpath.a_lt_b$in0[9] ;
 wire \dpath.a_lt_b$in1[0] ;
 wire \dpath.a_lt_b$in1[1] ;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net123;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net89;
 wire net107;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;

 BUFx4f_ASAP7_75t_R _297_ (.A(_029_),
    .Y(_084_));
 INVx1_ASAP7_75t_R _298_ (.A(_084_),
    .Y(_085_));
 BUFx6f_ASAP7_75t_R _299_ (.A(_085_),
    .Y(_086_));
 BUFx4f_ASAP7_75t_R _300_ (.A(_086_),
    .Y(net36));
 INVx1_ASAP7_75t_R _301_ (.A(_294_),
    .Y(\dpath.a_lt_b$in1[1] ));
 INVx2_ASAP7_75t_R _302_ (.A(_030_),
    .Y(\dpath.a_lt_b$in1[0] ));
 OA211x2_ASAP7_75t_R _303_ (.A1(_018_),
    .A2(net69),
    .B(_017_),
    .C(_015_),
    .Y(_087_));
 AO21x1_ASAP7_75t_R _304_ (.A1(net83),
    .A2(net89),
    .B(net72),
    .Y(_088_));
 OA21x2_ASAP7_75t_R _305_ (.A1(_087_),
    .A2(_088_),
    .B(_014_),
    .Y(_089_));
 OR2x2_ASAP7_75t_R _306_ (.A(net79),
    .B(_089_),
    .Y(_090_));
 AOI21x1_ASAP7_75t_R _307_ (.A1(_012_),
    .A2(_090_),
    .B(net95),
    .Y(_091_));
 INVx1_ASAP7_75t_R _308_ (.A(_028_),
    .Y(_092_));
 OA21x2_ASAP7_75t_R _309_ (.A1(_092_),
    .A2(net70),
    .B(_025_),
    .Y(_093_));
 OR3x1_ASAP7_75t_R _310_ (.A(net60),
    .B(net67),
    .C(net74),
    .Y(_094_));
 OA21x2_ASAP7_75t_R _311_ (.A1(net58),
    .A2(_023_),
    .B(_021_),
    .Y(_095_));
 OA21x2_ASAP7_75t_R _312_ (.A1(net76),
    .A2(_095_),
    .B(_020_),
    .Y(_096_));
 OA21x2_ASAP7_75t_R _313_ (.A1(_093_),
    .A2(_094_),
    .B(_096_),
    .Y(_097_));
 OR3x1_ASAP7_75t_R _314_ (.A(net69),
    .B(net61),
    .C(net56),
    .Y(_098_));
 NOR2x1_ASAP7_75t_R _315_ (.A(net78),
    .B(net73),
    .Y(_099_));
 INVx1_ASAP7_75t_R _316_ (.A(_099_),
    .Y(_100_));
 OR3x1_ASAP7_75t_R _317_ (.A(net93),
    .B(_098_),
    .C(_100_),
    .Y(_101_));
 OAI21x1_ASAP7_75t_R _318_ (.A1(_097_),
    .A2(net97),
    .B(_010_),
    .Y(_102_));
 OA21x2_ASAP7_75t_R _319_ (.A1(net114),
    .A2(net106),
    .B(_006_),
    .Y(_103_));
 OR2x2_ASAP7_75t_R _320_ (.A(_005_),
    .B(_103_),
    .Y(_104_));
 AO21x1_ASAP7_75t_R _321_ (.A1(_004_),
    .A2(_104_),
    .B(_047_),
    .Y(_105_));
 NAND2x1_ASAP7_75t_R _322_ (.A(_003_),
    .B(_105_),
    .Y(_106_));
 AO21x1_ASAP7_75t_R _323_ (.A1(net114),
    .A2(net92),
    .B(net105),
    .Y(_107_));
 AO21x1_ASAP7_75t_R _324_ (.A1(net112),
    .A2(_107_),
    .B(_005_),
    .Y(_108_));
 AO21x1_ASAP7_75t_R _325_ (.A1(_004_),
    .A2(_108_),
    .B(_047_),
    .Y(_109_));
 NAND2x1_ASAP7_75t_R _326_ (.A(_003_),
    .B(_109_),
    .Y(_110_));
 OA31x2_ASAP7_75t_R _327_ (.A1(_091_),
    .A2(_106_),
    .A3(_102_),
    .B1(_110_),
    .Y(_111_));
 BUFx4f_ASAP7_75t_R _328_ (.A(_111_),
    .Y(_112_));
 AND4x1_ASAP7_75t_R _329_ (.A(_286_),
    .B(_280_),
    .C(_281_),
    .D(_282_),
    .Y(_113_));
 AND5x1_ASAP7_75t_R _330_ (.A(_283_),
    .B(_284_),
    .C(_285_),
    .D(net101),
    .E(_113_),
    .Y(_114_));
 AND4x1_ASAP7_75t_R _331_ (.A(_287_),
    .B(_288_),
    .C(_289_),
    .D(_294_),
    .Y(_115_));
 AND4x1_ASAP7_75t_R _332_ (.A(_290_),
    .B(net98),
    .C(_292_),
    .D(net111),
    .Y(_116_));
 AND3x1_ASAP7_75t_R _333_ (.A(_114_),
    .B(_115_),
    .C(_116_),
    .Y(_117_));
 AO21x1_ASAP7_75t_R _334_ (.A1(_112_),
    .A2(_117_),
    .B(_045_),
    .Y(_118_));
 NAND2x1_ASAP7_75t_R _335_ (.A(net33),
    .B(net36),
    .Y(_119_));
 AOI21x1_ASAP7_75t_R _336_ (.A1(_118_),
    .A2(_119_),
    .B(net34),
    .Y(_002_));
 NAND2x1_ASAP7_75t_R _337_ (.A(_084_),
    .B(_045_),
    .Y(_120_));
 NOR2x1_ASAP7_75t_R _338_ (.A(_046_),
    .B(_120_),
    .Y(net53));
 INVx1_ASAP7_75t_R _339_ (.A(net33),
    .Y(_121_));
 BUFx6f_ASAP7_75t_R _340_ (.A(_085_),
    .Y(_122_));
 BUFx4f_ASAP7_75t_R _341_ (.A(_122_),
    .Y(_123_));
 AO221x1_ASAP7_75t_R _342_ (.A1(_121_),
    .A2(_123_),
    .B1(net53),
    .B2(net35),
    .C(net34),
    .Y(_000_));
 INVx2_ASAP7_75t_R _343_ (.A(_045_),
    .Y(_124_));
 AND3x1_ASAP7_75t_R _344_ (.A(_124_),
    .B(_112_),
    .C(_117_),
    .Y(_125_));
 AND2x6_ASAP7_75t_R _345_ (.A(_084_),
    .B(_045_),
    .Y(_126_));
 BUFx6f_ASAP7_75t_R _346_ (.A(_126_),
    .Y(_127_));
 AOI21x1_ASAP7_75t_R _347_ (.A1(net35),
    .A2(_127_),
    .B(_046_),
    .Y(_128_));
 INVx1_ASAP7_75t_R _348_ (.A(net34),
    .Y(_129_));
 OA21x2_ASAP7_75t_R _349_ (.A1(_125_),
    .A2(_128_),
    .B(_129_),
    .Y(_001_));
 INVx2_ASAP7_75t_R _350_ (.A(_031_),
    .Y(\dpath.a_lt_b$in0[9] ));
 INVx3_ASAP7_75t_R _351_ (.A(_032_),
    .Y(\dpath.a_lt_b$in0[8] ));
 INVx3_ASAP7_75t_R _352_ (.A(_033_),
    .Y(\dpath.a_lt_b$in0[7] ));
 INVx2_ASAP7_75t_R _353_ (.A(_034_),
    .Y(\dpath.a_lt_b$in0[6] ));
 INVx2_ASAP7_75t_R _354_ (.A(_035_),
    .Y(\dpath.a_lt_b$in0[5] ));
 INVx3_ASAP7_75t_R _355_ (.A(_036_),
    .Y(\dpath.a_lt_b$in0[4] ));
 INVx3_ASAP7_75t_R _356_ (.A(_037_),
    .Y(\dpath.a_lt_b$in0[3] ));
 INVx3_ASAP7_75t_R _357_ (.A(_038_),
    .Y(\dpath.a_lt_b$in0[2] ));
 INVx1_ASAP7_75t_R _358_ (.A(_279_),
    .Y(\dpath.a_lt_b$in0[1] ));
 INVx1_ASAP7_75t_R _359_ (.A(_039_),
    .Y(\dpath.a_lt_b$in0[15] ));
 INVx1_ASAP7_75t_R _360_ (.A(_040_),
    .Y(\dpath.a_lt_b$in0[14] ));
 INVx1_ASAP7_75t_R _361_ (.A(_041_),
    .Y(\dpath.a_lt_b$in0[13] ));
 INVx1_ASAP7_75t_R _362_ (.A(_042_),
    .Y(\dpath.a_lt_b$in0[12] ));
 INVx1_ASAP7_75t_R _363_ (.A(_043_),
    .Y(\dpath.a_lt_b$in0[11] ));
 INVx1_ASAP7_75t_R _364_ (.A(_044_),
    .Y(\dpath.a_lt_b$in0[10] ));
 AND2x4_ASAP7_75t_R _365_ (.A(_084_),
    .B(_124_),
    .Y(_130_));
 AND2x4_ASAP7_75t_R _366_ (.A(_111_),
    .B(_130_),
    .Y(_131_));
 NAND2x1_ASAP7_75t_R _367_ (.A(net37),
    .B(_131_),
    .Y(_132_));
 AO21x2_ASAP7_75t_R _368_ (.A1(_012_),
    .A2(_090_),
    .B(net94),
    .Y(_133_));
 OA21x2_ASAP7_75t_R _369_ (.A1(_101_),
    .A2(_097_),
    .B(_010_),
    .Y(_134_));
 AND3x4_ASAP7_75t_R _370_ (.A(_133_),
    .B(_134_),
    .C(_105_),
    .Y(_135_));
 AND3x1_ASAP7_75t_R _371_ (.A(_003_),
    .B(_084_),
    .C(_124_),
    .Y(_136_));
 OAI21x1_ASAP7_75t_R _372_ (.A1(_109_),
    .A2(_135_),
    .B(_136_),
    .Y(_137_));
 BUFx6f_ASAP7_75t_R _373_ (.A(net120),
    .Y(_138_));
 NAND2x1_ASAP7_75t_R _374_ (.A(_086_),
    .B(net8),
    .Y(_139_));
 OA211x2_ASAP7_75t_R _375_ (.A1(_030_),
    .A2(net119),
    .B(_139_),
    .C(_120_),
    .Y(_140_));
 AOI22x1_ASAP7_75t_R _376_ (.A1(_296_),
    .A2(_127_),
    .B1(_132_),
    .B2(_140_),
    .Y(_052_));
 BUFx4f_ASAP7_75t_R _377_ (.A(_124_),
    .Y(_141_));
 BUFx12f_ASAP7_75t_R _378_ (.A(net120),
    .Y(_142_));
 NOR2x2_ASAP7_75t_R _379_ (.A(_285_),
    .B(_142_),
    .Y(_143_));
 BUFx4f_ASAP7_75t_R _380_ (.A(_122_),
    .Y(_144_));
 AO21x1_ASAP7_75t_R _381_ (.A1(_144_),
    .A2(net19),
    .B(_127_),
    .Y(_145_));
 BUFx4f_ASAP7_75t_R _382_ (.A(_130_),
    .Y(_146_));
 OR2x2_ASAP7_75t_R _383_ (.A(net73),
    .B(_098_),
    .Y(_147_));
 OA21x2_ASAP7_75t_R _384_ (.A1(_097_),
    .A2(_147_),
    .B(_089_),
    .Y(_148_));
 XOR2x1_ASAP7_75t_R _385_ (.A(net77),
    .Y(net38),
    .B(_148_));
 AND3x1_ASAP7_75t_R _386_ (.A(_112_),
    .B(_146_),
    .C(net38),
    .Y(_149_));
 OA33x2_ASAP7_75t_R _387_ (.A1(net36),
    .A2(\dpath.a_lt_b$in0[10] ),
    .A3(_141_),
    .B1(_145_),
    .B2(_143_),
    .B3(_149_),
    .Y(_053_));
 NAND2x1_ASAP7_75t_R _388_ (.A(_086_),
    .B(net20),
    .Y(_150_));
 OA211x2_ASAP7_75t_R _389_ (.A1(_284_),
    .A2(net118),
    .B(_150_),
    .C(_120_),
    .Y(_151_));
 OA21x2_ASAP7_75t_R _390_ (.A1(net78),
    .A2(_014_),
    .B(_012_),
    .Y(_152_));
 INVx1_ASAP7_75t_R _391_ (.A(_295_),
    .Y(_278_));
 OA21x2_ASAP7_75t_R _392_ (.A1(_278_),
    .A2(_051_),
    .B(_027_),
    .Y(_153_));
 OR3x1_ASAP7_75t_R _393_ (.A(net80),
    .B(net65),
    .C(net58),
    .Y(_154_));
 OR3x1_ASAP7_75t_R _394_ (.A(_025_),
    .B(net58),
    .C(net65),
    .Y(_155_));
 OA211x2_ASAP7_75t_R _395_ (.A1(_153_),
    .A2(_154_),
    .B(_155_),
    .C(_095_),
    .Y(_156_));
 OR2x2_ASAP7_75t_R _396_ (.A(_098_),
    .B(net76),
    .Y(_157_));
 OR2x2_ASAP7_75t_R _397_ (.A(net62),
    .B(_020_),
    .Y(_158_));
 OR2x2_ASAP7_75t_R _398_ (.A(net56),
    .B(net69),
    .Y(_159_));
 AO21x1_ASAP7_75t_R _399_ (.A1(net81),
    .A2(_158_),
    .B(_159_),
    .Y(_160_));
 OA21x2_ASAP7_75t_R _400_ (.A1(_156_),
    .A2(_157_),
    .B(_160_),
    .Y(_161_));
 OA21x2_ASAP7_75t_R _401_ (.A1(net55),
    .A2(_017_),
    .B(net83),
    .Y(_162_));
 AO21x2_ASAP7_75t_R _402_ (.A1(_161_),
    .A2(_162_),
    .B(_100_),
    .Y(_163_));
 INVx1_ASAP7_75t_R _403_ (.A(net96),
    .Y(_164_));
 AO21x1_ASAP7_75t_R _404_ (.A1(_152_),
    .A2(net86),
    .B(_164_),
    .Y(_165_));
 NAND3x1_ASAP7_75t_R _405_ (.A(_164_),
    .B(_152_),
    .C(net86),
    .Y(_166_));
 NAND2x1_ASAP7_75t_R _406_ (.A(_112_),
    .B(_146_),
    .Y(_167_));
 AO21x1_ASAP7_75t_R _407_ (.A1(_165_),
    .A2(_166_),
    .B(_167_),
    .Y(_168_));
 AOI22x1_ASAP7_75t_R _408_ (.A1(_043_),
    .A2(_127_),
    .B1(_151_),
    .B2(_168_),
    .Y(_054_));
 OR2x2_ASAP7_75t_R _409_ (.A(_084_),
    .B(net21),
    .Y(_169_));
 NAND2x1_ASAP7_75t_R _410_ (.A(_042_),
    .B(_127_),
    .Y(_170_));
 OAI21x1_ASAP7_75t_R _411_ (.A1(_283_),
    .A2(_112_),
    .B(_146_),
    .Y(_171_));
 NAND2x2_ASAP7_75t_R _412_ (.A(_133_),
    .B(net122),
    .Y(_172_));
 XNOR2x1_ASAP7_75t_R _413_ (.B(_172_),
    .Y(net40),
    .A(net90));
 AO32x1_ASAP7_75t_R _414_ (.A1(_169_),
    .A2(_170_),
    .A3(_171_),
    .B1(net40),
    .B2(_131_),
    .Y(_055_));
 OA21x2_ASAP7_75t_R _415_ (.A1(net91),
    .A2(_010_),
    .B(_008_),
    .Y(_173_));
 AO21x1_ASAP7_75t_R _416_ (.A1(net93),
    .A2(_010_),
    .B(net91),
    .Y(_174_));
 AO32x1_ASAP7_75t_R _417_ (.A1(_152_),
    .A2(_163_),
    .A3(_173_),
    .B1(_174_),
    .B2(_008_),
    .Y(_175_));
 XOR2x1_ASAP7_75t_R _418_ (.A(_175_),
    .Y(net41),
    .B(net104));
 BUFx4f_ASAP7_75t_R _419_ (.A(_122_),
    .Y(_176_));
 AOI21x1_ASAP7_75t_R _420_ (.A1(_176_),
    .A2(net22),
    .B(_126_),
    .Y(_177_));
 OAI21x1_ASAP7_75t_R _421_ (.A1(_282_),
    .A2(net118),
    .B(_177_),
    .Y(_178_));
 NAND2x1_ASAP7_75t_R _422_ (.A(_041_),
    .B(_127_),
    .Y(_179_));
 AO32x1_ASAP7_75t_R _423_ (.A1(_112_),
    .A2(_146_),
    .A3(net41),
    .B1(_178_),
    .B2(_179_),
    .Y(_056_));
 OR2x2_ASAP7_75t_R _424_ (.A(_084_),
    .B(net24),
    .Y(_180_));
 NAND2x1_ASAP7_75t_R _425_ (.A(_040_),
    .B(_127_),
    .Y(_181_));
 OAI21x1_ASAP7_75t_R _426_ (.A1(_281_),
    .A2(_112_),
    .B(_146_),
    .Y(_182_));
 AO32x1_ASAP7_75t_R _427_ (.A1(_133_),
    .A2(_134_),
    .A3(_103_),
    .B1(_107_),
    .B2(net112),
    .Y(_183_));
 XOR2x1_ASAP7_75t_R _428_ (.A(_005_),
    .Y(net42),
    .B(_183_));
 AO32x1_ASAP7_75t_R _429_ (.A1(_180_),
    .A2(_181_),
    .A3(_182_),
    .B1(net42),
    .B2(_131_),
    .Y(_057_));
 OA21x2_ASAP7_75t_R _430_ (.A1(net105),
    .A2(_173_),
    .B(_006_),
    .Y(_184_));
 OA21x2_ASAP7_75t_R _431_ (.A1(_005_),
    .A2(_184_),
    .B(_152_),
    .Y(_185_));
 AND3x1_ASAP7_75t_R _432_ (.A(_185_),
    .B(_162_),
    .C(_161_),
    .Y(_186_));
 AO21x1_ASAP7_75t_R _433_ (.A1(net113),
    .A2(_174_),
    .B(net105),
    .Y(_187_));
 AND2x2_ASAP7_75t_R _434_ (.A(_100_),
    .B(_152_),
    .Y(_188_));
 AO221x1_ASAP7_75t_R _435_ (.A1(_006_),
    .A2(_187_),
    .B1(_188_),
    .B2(_184_),
    .C(_005_),
    .Y(_189_));
 OA21x2_ASAP7_75t_R _436_ (.A1(_186_),
    .A2(_189_),
    .B(_004_),
    .Y(_190_));
 XOR2x1_ASAP7_75t_R _437_ (.A(_047_),
    .Y(net43),
    .B(_190_));
 NAND2x1_ASAP7_75t_R _438_ (.A(_039_),
    .B(_126_),
    .Y(_191_));
 OAI21x1_ASAP7_75t_R _439_ (.A1(_280_),
    .A2(net117),
    .B(_130_),
    .Y(_192_));
 OA211x2_ASAP7_75t_R _440_ (.A1(_084_),
    .A2(net25),
    .B(_191_),
    .C(_192_),
    .Y(_193_));
 AO21x1_ASAP7_75t_R _441_ (.A1(_131_),
    .A2(net43),
    .B(_193_),
    .Y(_058_));
 AND3x1_ASAP7_75t_R _442_ (.A(net44),
    .B(_111_),
    .C(_130_),
    .Y(_194_));
 AO21x1_ASAP7_75t_R _443_ (.A1(_176_),
    .A2(net9),
    .B(_127_),
    .Y(_195_));
 BUFx12f_ASAP7_75t_R _444_ (.A(net120),
    .Y(_196_));
 NOR2x2_ASAP7_75t_R _445_ (.A(_294_),
    .B(_196_),
    .Y(_197_));
 OA33x2_ASAP7_75t_R _446_ (.A1(net36),
    .A2(\dpath.a_lt_b$in0[1] ),
    .A3(_141_),
    .B1(_194_),
    .B2(_195_),
    .B3(_197_),
    .Y(_059_));
 XNOR2x1_ASAP7_75t_R _447_ (.B(_028_),
    .Y(net45),
    .A(net71));
 AND3x1_ASAP7_75t_R _448_ (.A(_112_),
    .B(_146_),
    .C(net45),
    .Y(_198_));
 AO21x1_ASAP7_75t_R _449_ (.A1(_176_),
    .A2(net10),
    .B(_127_),
    .Y(_199_));
 NOR2x1_ASAP7_75t_R _450_ (.A(_293_),
    .B(_196_),
    .Y(_200_));
 OA33x2_ASAP7_75t_R _451_ (.A1(net36),
    .A2(net100),
    .A3(_141_),
    .B1(_198_),
    .B2(_199_),
    .B3(_200_),
    .Y(_060_));
 OA21x2_ASAP7_75t_R _452_ (.A1(net80),
    .A2(_153_),
    .B(_025_),
    .Y(_201_));
 XOR2x1_ASAP7_75t_R _453_ (.A(net66),
    .Y(net46),
    .B(_201_));
 AND3x1_ASAP7_75t_R _454_ (.A(_112_),
    .B(_146_),
    .C(net46),
    .Y(_202_));
 AO21x1_ASAP7_75t_R _455_ (.A1(_176_),
    .A2(net11),
    .B(_127_),
    .Y(_203_));
 NOR2x1_ASAP7_75t_R _456_ (.A(_292_),
    .B(_142_),
    .Y(_204_));
 OA33x2_ASAP7_75t_R _457_ (.A1(net36),
    .A2(\dpath.a_lt_b$in0[3] ),
    .A3(_141_),
    .B1(_202_),
    .B2(_203_),
    .B3(_204_),
    .Y(_061_));
 OA21x2_ASAP7_75t_R _458_ (.A1(net67),
    .A2(_093_),
    .B(net84),
    .Y(_205_));
 XOR2x1_ASAP7_75t_R _459_ (.A(net59),
    .Y(net47),
    .B(_205_));
 AND3x1_ASAP7_75t_R _460_ (.A(net117),
    .B(_146_),
    .C(net47),
    .Y(_206_));
 AO21x1_ASAP7_75t_R _461_ (.A1(_176_),
    .A2(net13),
    .B(_126_),
    .Y(_207_));
 NOR2x1_ASAP7_75t_R _462_ (.A(net99),
    .B(_142_),
    .Y(_208_));
 OA33x2_ASAP7_75t_R _463_ (.A1(net36),
    .A2(net87),
    .A3(_141_),
    .B1(_206_),
    .B2(_207_),
    .B3(_208_),
    .Y(_062_));
 XOR2x1_ASAP7_75t_R _464_ (.A(net75),
    .Y(net48),
    .B(net85));
 AND3x1_ASAP7_75t_R _465_ (.A(net117),
    .B(_146_),
    .C(net48),
    .Y(_209_));
 AO21x1_ASAP7_75t_R _466_ (.A1(_176_),
    .A2(net14),
    .B(_126_),
    .Y(_210_));
 NOR2x1_ASAP7_75t_R _467_ (.A(_290_),
    .B(net118),
    .Y(_211_));
 OA33x2_ASAP7_75t_R _468_ (.A1(net36),
    .A2(\dpath.a_lt_b$in0[5] ),
    .A3(_141_),
    .B1(_209_),
    .B2(_210_),
    .B3(_211_),
    .Y(_063_));
 XOR2x1_ASAP7_75t_R _469_ (.A(net102),
    .Y(net49),
    .B(net63));
 AND3x1_ASAP7_75t_R _470_ (.A(net117),
    .B(_130_),
    .C(net49),
    .Y(_212_));
 AO21x1_ASAP7_75t_R _471_ (.A1(_176_),
    .A2(net15),
    .B(_126_),
    .Y(_213_));
 NOR2x1_ASAP7_75t_R _472_ (.A(_289_),
    .B(net118),
    .Y(_214_));
 OA33x2_ASAP7_75t_R _473_ (.A1(net36),
    .A2(\dpath.a_lt_b$in0[6] ),
    .A3(_141_),
    .B1(_212_),
    .B2(_213_),
    .B3(_214_),
    .Y(_064_));
 OR3x1_ASAP7_75t_R _474_ (.A(net64),
    .B(net76),
    .C(_156_),
    .Y(_215_));
 AND3x1_ASAP7_75t_R _475_ (.A(_215_),
    .B(_158_),
    .C(net82),
    .Y(_216_));
 XOR2x1_ASAP7_75t_R _476_ (.A(net68),
    .Y(net50),
    .B(_216_));
 AND2x2_ASAP7_75t_R _477_ (.A(_131_),
    .B(net50),
    .Y(_217_));
 AO21x1_ASAP7_75t_R _478_ (.A1(_176_),
    .A2(net16),
    .B(_126_),
    .Y(_218_));
 NOR2x1_ASAP7_75t_R _479_ (.A(_288_),
    .B(_142_),
    .Y(_219_));
 OA33x2_ASAP7_75t_R _480_ (.A1(net36),
    .A2(\dpath.a_lt_b$in0[7] ),
    .A3(_141_),
    .B1(_217_),
    .B2(_218_),
    .B3(_219_),
    .Y(_065_));
 NOR2x1_ASAP7_75t_R _481_ (.A(_287_),
    .B(net118),
    .Y(_220_));
 AO21x1_ASAP7_75t_R _482_ (.A1(_176_),
    .A2(net17),
    .B(_126_),
    .Y(_221_));
 OA21x2_ASAP7_75t_R _483_ (.A1(_097_),
    .A2(net61),
    .B(_018_),
    .Y(_222_));
 OA21x2_ASAP7_75t_R _484_ (.A1(net69),
    .A2(_222_),
    .B(_017_),
    .Y(_223_));
 XOR2x1_ASAP7_75t_R _485_ (.A(net57),
    .Y(net51),
    .B(_223_));
 AND3x1_ASAP7_75t_R _486_ (.A(_112_),
    .B(_146_),
    .C(net51),
    .Y(_224_));
 OA33x2_ASAP7_75t_R _487_ (.A1(_123_),
    .A2(\dpath.a_lt_b$in0[8] ),
    .A3(_141_),
    .B1(_220_),
    .B2(_221_),
    .B3(_224_),
    .Y(_066_));
 NOR2x1_ASAP7_75t_R _488_ (.A(_286_),
    .B(_142_),
    .Y(_225_));
 AO21x1_ASAP7_75t_R _489_ (.A1(_176_),
    .A2(net18),
    .B(_126_),
    .Y(_226_));
 NAND2x1_ASAP7_75t_R _490_ (.A(_161_),
    .B(_162_),
    .Y(_227_));
 XNOR2x1_ASAP7_75t_R _491_ (.B(_227_),
    .Y(net52),
    .A(net72));
 AND2x2_ASAP7_75t_R _492_ (.A(_131_),
    .B(net52),
    .Y(_228_));
 OA33x2_ASAP7_75t_R _493_ (.A1(_123_),
    .A2(\dpath.a_lt_b$in0[9] ),
    .A3(_141_),
    .B1(_225_),
    .B2(_226_),
    .B3(_228_),
    .Y(_067_));
 BUFx12f_ASAP7_75t_R _494_ (.A(net120),
    .Y(_229_));
 AND2x2_ASAP7_75t_R _495_ (.A(_084_),
    .B(\dpath.a_lt_b$in1[0] ),
    .Y(_230_));
 AO21x1_ASAP7_75t_R _496_ (.A1(_123_),
    .A2(net1),
    .B(_230_),
    .Y(_231_));
 NOR2x1_ASAP7_75t_R _497_ (.A(net103),
    .B(net116),
    .Y(_232_));
 AO21x1_ASAP7_75t_R _498_ (.A1(net123),
    .A2(_231_),
    .B(_232_),
    .Y(_068_));
 NOR2x1_ASAP7_75t_R _499_ (.A(\dpath.a_lt_b$in0[10] ),
    .B(_229_),
    .Y(_233_));
 NAND2x1_ASAP7_75t_R _500_ (.A(_086_),
    .B(net2),
    .Y(_234_));
 OA211x2_ASAP7_75t_R _501_ (.A1(_123_),
    .A2(_285_),
    .B(_138_),
    .C(_234_),
    .Y(_235_));
 NOR2x1_ASAP7_75t_R _502_ (.A(_233_),
    .B(_235_),
    .Y(_069_));
 NOR2x1_ASAP7_75t_R _503_ (.A(\dpath.a_lt_b$in0[11] ),
    .B(_229_),
    .Y(_236_));
 NAND2x1_ASAP7_75t_R _504_ (.A(_086_),
    .B(net3),
    .Y(_237_));
 OA211x2_ASAP7_75t_R _505_ (.A1(_123_),
    .A2(_284_),
    .B(_138_),
    .C(_237_),
    .Y(_238_));
 NOR2x1_ASAP7_75t_R _506_ (.A(_236_),
    .B(_238_),
    .Y(_070_));
 NOR2x1_ASAP7_75t_R _507_ (.A(\dpath.a_lt_b$in0[12] ),
    .B(_229_),
    .Y(_239_));
 NAND2x1_ASAP7_75t_R _508_ (.A(_086_),
    .B(net4),
    .Y(_240_));
 OA211x2_ASAP7_75t_R _509_ (.A1(_123_),
    .A2(_283_),
    .B(_138_),
    .C(_240_),
    .Y(_241_));
 NOR2x1_ASAP7_75t_R _510_ (.A(_239_),
    .B(_241_),
    .Y(_071_));
 NOR2x1_ASAP7_75t_R _511_ (.A(\dpath.a_lt_b$in0[13] ),
    .B(_229_),
    .Y(_242_));
 NAND2x1_ASAP7_75t_R _512_ (.A(_086_),
    .B(net5),
    .Y(_243_));
 OA211x2_ASAP7_75t_R _513_ (.A1(_123_),
    .A2(_282_),
    .B(_138_),
    .C(_243_),
    .Y(_244_));
 NOR2x1_ASAP7_75t_R _514_ (.A(_242_),
    .B(_244_),
    .Y(_072_));
 NOR2x1_ASAP7_75t_R _515_ (.A(\dpath.a_lt_b$in0[14] ),
    .B(_229_),
    .Y(_245_));
 NAND2x1_ASAP7_75t_R _516_ (.A(_086_),
    .B(net6),
    .Y(_246_));
 OA211x2_ASAP7_75t_R _517_ (.A1(_123_),
    .A2(_281_),
    .B(_138_),
    .C(_246_),
    .Y(_247_));
 NOR2x1_ASAP7_75t_R _518_ (.A(_245_),
    .B(_247_),
    .Y(_073_));
 NOR2x1_ASAP7_75t_R _519_ (.A(\dpath.a_lt_b$in0[15] ),
    .B(net123),
    .Y(_248_));
 NAND2x1_ASAP7_75t_R _520_ (.A(_086_),
    .B(net7),
    .Y(_249_));
 OA211x2_ASAP7_75t_R _521_ (.A1(_144_),
    .A2(_280_),
    .B(net119),
    .C(_249_),
    .Y(_250_));
 NOR2x1_ASAP7_75t_R _522_ (.A(_248_),
    .B(_250_),
    .Y(_074_));
 AND2x2_ASAP7_75t_R _523_ (.A(_084_),
    .B(\dpath.a_lt_b$in1[1] ),
    .Y(_251_));
 AO21x1_ASAP7_75t_R _524_ (.A1(_123_),
    .A2(net12),
    .B(_251_),
    .Y(_252_));
 NOR2x1_ASAP7_75t_R _525_ (.A(_279_),
    .B(net116),
    .Y(_253_));
 AO21x1_ASAP7_75t_R _526_ (.A1(net123),
    .A2(_252_),
    .B(_253_),
    .Y(_075_));
 NOR2x1_ASAP7_75t_R _527_ (.A(net100),
    .B(net123),
    .Y(_254_));
 NAND2x1_ASAP7_75t_R _528_ (.A(_086_),
    .B(net23),
    .Y(_255_));
 OA211x2_ASAP7_75t_R _529_ (.A1(_144_),
    .A2(_293_),
    .B(net119),
    .C(_255_),
    .Y(_256_));
 NOR2x1_ASAP7_75t_R _530_ (.A(_254_),
    .B(_256_),
    .Y(_076_));
 NOR2x1_ASAP7_75t_R _531_ (.A(\dpath.a_lt_b$in0[3] ),
    .B(net123),
    .Y(_257_));
 NAND2x1_ASAP7_75t_R _532_ (.A(_122_),
    .B(net26),
    .Y(_258_));
 OA211x2_ASAP7_75t_R _533_ (.A1(_144_),
    .A2(_292_),
    .B(net119),
    .C(_258_),
    .Y(_259_));
 NOR2x1_ASAP7_75t_R _534_ (.A(_257_),
    .B(_259_),
    .Y(_077_));
 NOR2x2_ASAP7_75t_R _535_ (.A(net87),
    .B(_196_),
    .Y(_260_));
 NAND2x1_ASAP7_75t_R _536_ (.A(_122_),
    .B(net27),
    .Y(_261_));
 OA211x2_ASAP7_75t_R _537_ (.A1(_144_),
    .A2(_291_),
    .B(net119),
    .C(_261_),
    .Y(_262_));
 NOR2x1_ASAP7_75t_R _538_ (.A(_262_),
    .B(_260_),
    .Y(_078_));
 NOR2x1_ASAP7_75t_R _539_ (.A(\dpath.a_lt_b$in0[5] ),
    .B(_196_),
    .Y(_263_));
 NAND2x1_ASAP7_75t_R _540_ (.A(_122_),
    .B(net28),
    .Y(_264_));
 OA211x2_ASAP7_75t_R _541_ (.A1(_144_),
    .A2(_290_),
    .B(net115),
    .C(_264_),
    .Y(_265_));
 NOR2x1_ASAP7_75t_R _542_ (.A(_263_),
    .B(_265_),
    .Y(_079_));
 NOR2x1_ASAP7_75t_R _543_ (.A(\dpath.a_lt_b$in0[6] ),
    .B(net116),
    .Y(_266_));
 NAND2x1_ASAP7_75t_R _544_ (.A(_122_),
    .B(net29),
    .Y(_267_));
 OA211x2_ASAP7_75t_R _545_ (.A1(_144_),
    .A2(_289_),
    .B(net115),
    .C(_267_),
    .Y(_268_));
 NOR2x1_ASAP7_75t_R _546_ (.A(_266_),
    .B(_268_),
    .Y(_080_));
 NOR2x1_ASAP7_75t_R _547_ (.A(net88),
    .B(net116),
    .Y(_269_));
 NAND2x1_ASAP7_75t_R _548_ (.A(_122_),
    .B(net30),
    .Y(_270_));
 OA211x2_ASAP7_75t_R _549_ (.A1(_144_),
    .A2(_288_),
    .B(net115),
    .C(_270_),
    .Y(_271_));
 NOR2x1_ASAP7_75t_R _550_ (.A(_269_),
    .B(_271_),
    .Y(_081_));
 NOR2x1_ASAP7_75t_R _551_ (.A(net121),
    .B(net116),
    .Y(_272_));
 NAND2x1_ASAP7_75t_R _552_ (.A(_122_),
    .B(net31),
    .Y(_273_));
 OA211x2_ASAP7_75t_R _553_ (.A1(_144_),
    .A2(_287_),
    .B(net115),
    .C(_273_),
    .Y(_274_));
 NOR2x1_ASAP7_75t_R _554_ (.A(_272_),
    .B(_274_),
    .Y(_082_));
 NOR2x1_ASAP7_75t_R _555_ (.A(\dpath.a_lt_b$in0[9] ),
    .B(_196_),
    .Y(_275_));
 NAND2x1_ASAP7_75t_R _556_ (.A(_122_),
    .B(net32),
    .Y(_276_));
 OA211x2_ASAP7_75t_R _557_ (.A1(_144_),
    .A2(_286_),
    .B(_137_),
    .C(_276_),
    .Y(_277_));
 NOR2x1_ASAP7_75t_R _558_ (.A(_275_),
    .B(_277_),
    .Y(_083_));
 NAND2x1_ASAP7_75t_R _559_ (.A(_166_),
    .B(_165_),
    .Y(net39));
 FAx1_ASAP7_75t_R _560_ (.SN(net44),
    .A(_279_),
    .B(\dpath.a_lt_b$in1[1] ),
    .CI(_278_),
    .CON(_028_));
 HAxp5_ASAP7_75t_R _561_ (.A(_280_),
    .B(\dpath.a_lt_b$in0[15] ),
    .CON(_003_),
    .SN(_047_));
 HAxp5_ASAP7_75t_R _562_ (.A(_281_),
    .B(\dpath.a_lt_b$in0[14] ),
    .CON(_004_),
    .SN(_005_));
 HAxp5_ASAP7_75t_R _563_ (.A(\dpath.a_lt_b$in0[13] ),
    .B(_282_),
    .CON(_006_),
    .SN(_007_));
 HAxp5_ASAP7_75t_R _564_ (.A(\dpath.a_lt_b$in0[12] ),
    .B(_283_),
    .CON(_008_),
    .SN(_009_));
 HAxp5_ASAP7_75t_R _565_ (.A(\dpath.a_lt_b$in0[11] ),
    .B(_284_),
    .CON(_010_),
    .SN(_011_));
 HAxp5_ASAP7_75t_R _566_ (.A(\dpath.a_lt_b$in0[10] ),
    .B(_285_),
    .CON(_012_),
    .SN(_013_));
 HAxp5_ASAP7_75t_R _567_ (.A(\dpath.a_lt_b$in0[9] ),
    .B(_286_),
    .CON(_014_),
    .SN(_048_));
 HAxp5_ASAP7_75t_R _568_ (.A(_287_),
    .B(\dpath.a_lt_b$in0[8] ),
    .CON(_015_),
    .SN(_016_));
 HAxp5_ASAP7_75t_R _569_ (.A(\dpath.a_lt_b$in0[7] ),
    .B(_288_),
    .CON(_017_),
    .SN(_049_));
 HAxp5_ASAP7_75t_R _570_ (.A(\dpath.a_lt_b$in0[6] ),
    .B(_289_),
    .CON(_018_),
    .SN(_019_));
 HAxp5_ASAP7_75t_R _571_ (.A(\dpath.a_lt_b$in0[5] ),
    .B(_290_),
    .CON(_020_),
    .SN(_050_));
 HAxp5_ASAP7_75t_R _572_ (.A(\dpath.a_lt_b$in0[4] ),
    .B(_291_),
    .CON(_021_),
    .SN(_022_));
 HAxp5_ASAP7_75t_R _573_ (.A(\dpath.a_lt_b$in0[3] ),
    .B(_292_),
    .CON(_023_),
    .SN(_024_));
 HAxp5_ASAP7_75t_R _574_ (.A(_293_),
    .B(\dpath.a_lt_b$in0[2] ),
    .CON(_025_),
    .SN(_026_));
 HAxp5_ASAP7_75t_R _575_ (.A(_294_),
    .B(\dpath.a_lt_b$in0[1] ),
    .CON(_027_),
    .SN(_051_));
 HAxp5_ASAP7_75t_R _576_ (.A(\dpath.a_lt_b$in1[0] ),
    .B(_296_),
    .CON(_295_),
    .SN(net37));
 DFFHQNx1_ASAP7_75t_R \ctrl.state.out[0]$_DFF_P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_000_),
    .QN(_029_));
 DFFHQNx2_ASAP7_75t_R \ctrl.state.out[1]$_DFF_P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_001_),
    .QN(_046_));
 DFFHQNx2_ASAP7_75t_R \ctrl.state.out[2]$_DFF_P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_002_),
    .QN(_045_));
 DFFHQNx2_ASAP7_75t_R \dpath.a_reg.out[0]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .D(_052_),
    .QN(_296_));
 DFFHQNx3_ASAP7_75t_R \dpath.a_reg.out[10]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .D(_053_),
    .QN(_044_));
 DFFHQNx2_ASAP7_75t_R \dpath.a_reg.out[11]$_DFFE_PP_  (.CLK(clknet_2_3__leaf_clk),
    .D(_054_),
    .QN(_043_));
 DFFHQNx2_ASAP7_75t_R \dpath.a_reg.out[12]$_DFFE_PP_  (.CLK(clknet_2_3__leaf_clk),
    .D(_055_),
    .QN(_042_));
 DFFHQNx2_ASAP7_75t_R \dpath.a_reg.out[13]$_DFFE_PP_  (.CLK(clknet_2_2__leaf_clk),
    .D(_056_),
    .QN(_041_));
 DFFHQNx2_ASAP7_75t_R \dpath.a_reg.out[14]$_DFFE_PP_  (.CLK(clknet_2_2__leaf_clk),
    .D(_057_),
    .QN(_040_));
 DFFHQNx2_ASAP7_75t_R \dpath.a_reg.out[15]$_DFFE_PP_  (.CLK(clknet_2_2__leaf_clk),
    .D(_058_),
    .QN(_039_));
 DFFHQNx2_ASAP7_75t_R \dpath.a_reg.out[1]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .D(_059_),
    .QN(_279_));
 DFFHQNx3_ASAP7_75t_R \dpath.a_reg.out[2]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .D(_060_),
    .QN(_038_));
 DFFHQNx3_ASAP7_75t_R \dpath.a_reg.out[3]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .D(_061_),
    .QN(_037_));
 DFFHQNx3_ASAP7_75t_R \dpath.a_reg.out[4]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .D(_062_),
    .QN(_036_));
 DFFHQNx3_ASAP7_75t_R \dpath.a_reg.out[5]$_DFFE_PP_  (.CLK(clknet_2_0__leaf_clk),
    .D(_063_),
    .QN(_035_));
 DFFHQNx3_ASAP7_75t_R \dpath.a_reg.out[6]$_DFFE_PP_  (.CLK(clknet_2_0__leaf_clk),
    .D(_064_),
    .QN(_034_));
 DFFHQNx3_ASAP7_75t_R \dpath.a_reg.out[7]$_DFFE_PP_  (.CLK(clknet_2_0__leaf_clk),
    .D(_065_),
    .QN(_033_));
 DFFHQNx3_ASAP7_75t_R \dpath.a_reg.out[8]$_DFFE_PP_  (.CLK(clknet_2_0__leaf_clk),
    .D(_066_),
    .QN(_032_));
 DFFHQNx3_ASAP7_75t_R \dpath.a_reg.out[9]$_DFFE_PP_  (.CLK(clknet_2_2__leaf_clk),
    .D(_067_),
    .QN(_031_));
 DFFHQNx2_ASAP7_75t_R \dpath.b_reg.out[0]$_DFFE_PP_  (.CLK(clknet_2_3__leaf_clk),
    .D(_068_),
    .QN(_030_));
 DFFHQNx2_ASAP7_75t_R \dpath.b_reg.out[10]$_DFFE_PP_  (.CLK(clknet_2_3__leaf_clk),
    .D(_069_),
    .QN(_285_));
 DFFHQNx2_ASAP7_75t_R \dpath.b_reg.out[11]$_DFFE_PP_  (.CLK(clknet_2_3__leaf_clk),
    .D(_070_),
    .QN(_284_));
 DFFHQNx2_ASAP7_75t_R \dpath.b_reg.out[12]$_DFFE_PP_  (.CLK(clknet_2_3__leaf_clk),
    .D(_071_),
    .QN(_283_));
 DFFHQNx2_ASAP7_75t_R \dpath.b_reg.out[13]$_DFFE_PP_  (.CLK(clknet_2_2__leaf_clk),
    .D(_072_),
    .QN(_282_));
 DFFHQNx2_ASAP7_75t_R \dpath.b_reg.out[14]$_DFFE_PP_  (.CLK(clknet_2_2__leaf_clk),
    .D(_073_),
    .QN(_281_));
 DFFHQNx2_ASAP7_75t_R \dpath.b_reg.out[15]$_DFFE_PP_  (.CLK(clknet_2_2__leaf_clk),
    .D(_074_),
    .QN(_280_));
 DFFHQNx2_ASAP7_75t_R \dpath.b_reg.out[1]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .D(_075_),
    .QN(_294_));
 DFFHQNx2_ASAP7_75t_R \dpath.b_reg.out[2]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .D(_076_),
    .QN(_293_));
 DFFHQNx2_ASAP7_75t_R \dpath.b_reg.out[3]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .D(_077_),
    .QN(_292_));
 DFFHQNx2_ASAP7_75t_R \dpath.b_reg.out[4]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .D(_078_),
    .QN(_291_));
 DFFHQNx2_ASAP7_75t_R \dpath.b_reg.out[5]$_DFFE_PP_  (.CLK(clknet_2_0__leaf_clk),
    .D(_079_),
    .QN(_290_));
 DFFHQNx2_ASAP7_75t_R \dpath.b_reg.out[6]$_DFFE_PP_  (.CLK(clknet_2_0__leaf_clk),
    .D(_080_),
    .QN(_289_));
 DFFHQNx2_ASAP7_75t_R \dpath.b_reg.out[7]$_DFFE_PP_  (.CLK(clknet_2_0__leaf_clk),
    .D(_081_),
    .QN(_288_));
 DFFHQNx2_ASAP7_75t_R \dpath.b_reg.out[8]$_DFFE_PP_  (.CLK(clknet_2_0__leaf_clk),
    .D(_082_),
    .QN(_287_));
 DFFHQNx2_ASAP7_75t_R \dpath.b_reg.out[9]$_DFFE_PP_  (.CLK(clknet_2_2__leaf_clk),
    .D(_083_),
    .QN(_286_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Left_52 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Left_53 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Left_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Left_55 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Left_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Left_57 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Left_58 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Left_59 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Left_60 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Left_61 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Left_62 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Left_63 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Left_64 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Left_65 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Left_66 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Left_67 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Left_68 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Left_69 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Left_70 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Left_71 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Left_72 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Left_73 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Left_74 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Left_75 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Left_76 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Left_77 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Left_78 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Left_79 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Left_80 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Left_81 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Left_82 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Left_83 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Left_84 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Left_85 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Left_86 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Left_87 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Left_88 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Left_89 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Left_90 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Left_91 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Left_92 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Left_93 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Left_94 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Left_95 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Left_96 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Left_97 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Left_98 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Left_99 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Left_100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Left_101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Left_102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Left_103 ();
 BUFx2_ASAP7_75t_R input1 (.A(req_msg[0]),
    .Y(net1));
 BUFx2_ASAP7_75t_R input2 (.A(req_msg[10]),
    .Y(net2));
 BUFx2_ASAP7_75t_R input3 (.A(req_msg[11]),
    .Y(net3));
 BUFx2_ASAP7_75t_R input4 (.A(req_msg[12]),
    .Y(net4));
 BUFx2_ASAP7_75t_R input5 (.A(req_msg[13]),
    .Y(net5));
 BUFx2_ASAP7_75t_R input6 (.A(req_msg[14]),
    .Y(net6));
 BUFx2_ASAP7_75t_R input7 (.A(req_msg[15]),
    .Y(net7));
 BUFx2_ASAP7_75t_R input8 (.A(req_msg[16]),
    .Y(net8));
 BUFx2_ASAP7_75t_R input9 (.A(req_msg[17]),
    .Y(net9));
 BUFx2_ASAP7_75t_R input10 (.A(req_msg[18]),
    .Y(net10));
 BUFx2_ASAP7_75t_R input11 (.A(req_msg[19]),
    .Y(net11));
 BUFx2_ASAP7_75t_R input12 (.A(req_msg[1]),
    .Y(net12));
 BUFx2_ASAP7_75t_R input13 (.A(req_msg[20]),
    .Y(net13));
 BUFx2_ASAP7_75t_R input14 (.A(req_msg[21]),
    .Y(net14));
 BUFx2_ASAP7_75t_R input15 (.A(req_msg[22]),
    .Y(net15));
 BUFx2_ASAP7_75t_R input16 (.A(req_msg[23]),
    .Y(net16));
 BUFx2_ASAP7_75t_R input17 (.A(req_msg[24]),
    .Y(net17));
 BUFx2_ASAP7_75t_R input18 (.A(req_msg[25]),
    .Y(net18));
 BUFx2_ASAP7_75t_R input19 (.A(req_msg[26]),
    .Y(net19));
 BUFx2_ASAP7_75t_R input20 (.A(req_msg[27]),
    .Y(net20));
 BUFx2_ASAP7_75t_R input21 (.A(req_msg[28]),
    .Y(net21));
 BUFx2_ASAP7_75t_R input22 (.A(req_msg[29]),
    .Y(net22));
 BUFx2_ASAP7_75t_R input23 (.A(req_msg[2]),
    .Y(net23));
 BUFx2_ASAP7_75t_R input24 (.A(req_msg[30]),
    .Y(net24));
 BUFx2_ASAP7_75t_R input25 (.A(req_msg[31]),
    .Y(net25));
 BUFx2_ASAP7_75t_R input26 (.A(req_msg[3]),
    .Y(net26));
 BUFx2_ASAP7_75t_R input27 (.A(req_msg[4]),
    .Y(net27));
 BUFx2_ASAP7_75t_R input28 (.A(req_msg[5]),
    .Y(net28));
 BUFx2_ASAP7_75t_R input29 (.A(req_msg[6]),
    .Y(net29));
 BUFx2_ASAP7_75t_R input30 (.A(req_msg[7]),
    .Y(net30));
 BUFx2_ASAP7_75t_R input31 (.A(req_msg[8]),
    .Y(net31));
 BUFx2_ASAP7_75t_R input32 (.A(req_msg[9]),
    .Y(net32));
 BUFx2_ASAP7_75t_R input33 (.A(req_val),
    .Y(net33));
 BUFx2_ASAP7_75t_R input34 (.A(reset),
    .Y(net34));
 BUFx2_ASAP7_75t_R input35 (.A(resp_rdy),
    .Y(net35));
 BUFx2_ASAP7_75t_R output36 (.A(net36),
    .Y(req_rdy));
 BUFx2_ASAP7_75t_R output37 (.A(net37),
    .Y(resp_msg[0]));
 BUFx2_ASAP7_75t_R output38 (.A(net38),
    .Y(resp_msg[10]));
 BUFx2_ASAP7_75t_R output39 (.A(net39),
    .Y(resp_msg[11]));
 BUFx2_ASAP7_75t_R output40 (.A(net40),
    .Y(resp_msg[12]));
 BUFx3_ASAP7_75t_R output41 (.A(net41),
    .Y(resp_msg[13]));
 BUFx2_ASAP7_75t_R output42 (.A(net42),
    .Y(resp_msg[14]));
 BUFx2_ASAP7_75t_R output43 (.A(net43),
    .Y(resp_msg[15]));
 BUFx2_ASAP7_75t_R output44 (.A(net44),
    .Y(resp_msg[1]));
 BUFx2_ASAP7_75t_R output45 (.A(net45),
    .Y(resp_msg[2]));
 BUFx2_ASAP7_75t_R output46 (.A(net46),
    .Y(resp_msg[3]));
 BUFx2_ASAP7_75t_R output47 (.A(net47),
    .Y(resp_msg[4]));
 BUFx2_ASAP7_75t_R output48 (.A(net48),
    .Y(resp_msg[5]));
 BUFx3_ASAP7_75t_R output49 (.A(net49),
    .Y(resp_msg[6]));
 BUFx2_ASAP7_75t_R output50 (.A(net50),
    .Y(resp_msg[7]));
 BUFx2_ASAP7_75t_R output51 (.A(net51),
    .Y(resp_msg[8]));
 BUFx2_ASAP7_75t_R output52 (.A(net52),
    .Y(resp_msg[9]));
 BUFx2_ASAP7_75t_R output53 (.A(net53),
    .Y(resp_val));
 BUFx2_ASAP7_75t_R clkbuf_0_clk (.A(clk),
    .Y(clknet_0_clk));
 BUFx2_ASAP7_75t_R clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Y(clknet_2_0__leaf_clk));
 BUFx2_ASAP7_75t_R clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Y(clknet_2_1__leaf_clk));
 BUFx2_ASAP7_75t_R clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Y(clknet_2_2__leaf_clk));
 BUFx2_ASAP7_75t_R clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Y(clknet_2_3__leaf_clk));
 BUFx4f_ASAP7_75t_R clkload0 (.A(clknet_2_0__leaf_clk));
 BUFx4f_ASAP7_75t_R clkload1 (.A(clknet_2_2__leaf_clk));
 INVxp67_ASAP7_75t_R clkload2 (.A(clknet_2_3__leaf_clk));
 BUFx12f_ASAP7_75t_R clone70 (.A(net120),
    .Y(net123));
 BUFx2_ASAP7_75t_R rebuffer2 (.A(net89),
    .Y(net55));
 BUFx3_ASAP7_75t_R rebuffer3 (.A(_016_),
    .Y(net56));
 BUFx2_ASAP7_75t_R rebuffer4 (.A(net56),
    .Y(net57));
 BUFx3_ASAP7_75t_R rebuffer5 (.A(_022_),
    .Y(net58));
 BUFx2_ASAP7_75t_R rebuffer6 (.A(net58),
    .Y(net59));
 BUFx2_ASAP7_75t_R rebuffer7 (.A(_022_),
    .Y(net60));
 BUFx3_ASAP7_75t_R rebuffer8 (.A(_019_),
    .Y(net61));
 BUFx2_ASAP7_75t_R rebuffer9 (.A(net61),
    .Y(net62));
 BUFx2_ASAP7_75t_R rebuffer10 (.A(net62),
    .Y(net63));
 BUFx2_ASAP7_75t_R rebuffer11 (.A(net62),
    .Y(net64));
 BUFx3_ASAP7_75t_R rebuffer12 (.A(_024_),
    .Y(net65));
 BUFx2_ASAP7_75t_R rebuffer13 (.A(net65),
    .Y(net66));
 BUFx2_ASAP7_75t_R rebuffer14 (.A(net65),
    .Y(net67));
 BUFx2_ASAP7_75t_R rebuffer15 (.A(net107),
    .Y(net68));
 BUFx3_ASAP7_75t_R rebuffer16 (.A(_049_),
    .Y(net69));
 BUFx3_ASAP7_75t_R rebuffer17 (.A(net80),
    .Y(net70));
 BUFx2_ASAP7_75t_R rebuffer18 (.A(_026_),
    .Y(net71));
 BUFx3_ASAP7_75t_R rebuffer19 (.A(_048_),
    .Y(net72));
 BUFx2_ASAP7_75t_R rebuffer20 (.A(net72),
    .Y(net73));
 BUFx2_ASAP7_75t_R rebuffer21 (.A(_050_),
    .Y(net74));
 BUFx3_ASAP7_75t_R rebuffer22 (.A(_050_),
    .Y(net75));
 BUFx3_ASAP7_75t_R rebuffer23 (.A(net75),
    .Y(net76));
 BUFx2_ASAP7_75t_R rebuffer24 (.A(_013_),
    .Y(net77));
 BUFx3_ASAP7_75t_R rebuffer25 (.A(_013_),
    .Y(net78));
 BUFx2_ASAP7_75t_R rebuffer26 (.A(net78),
    .Y(net79));
 BUFx3_ASAP7_75t_R rebuffer27 (.A(_026_),
    .Y(net80));
 BUFx2_ASAP7_75t_R rebuffer28 (.A(_018_),
    .Y(net81));
 BUFx2_ASAP7_75t_R rebuffer29 (.A(net81),
    .Y(net82));
 BUFx3_ASAP7_75t_R rebuffer30 (.A(_015_),
    .Y(net83));
 BUFx2_ASAP7_75t_R rebuffer31 (.A(_023_),
    .Y(net84));
 BUFx2_ASAP7_75t_R rebuffer32 (.A(_156_),
    .Y(net85));
 BUFx2_ASAP7_75t_R rebuffer33 (.A(_163_),
    .Y(net86));
 BUFx2_ASAP7_75t_R rebuffer34 (.A(\dpath.a_lt_b$in0[4] ),
    .Y(net87));
 BUFx2_ASAP7_75t_R rebuffer35 (.A(\dpath.a_lt_b$in0[7] ),
    .Y(net88));
 BUFx2_ASAP7_75t_R rebuffer37 (.A(_009_),
    .Y(net90));
 BUFx3_ASAP7_75t_R rebuffer38 (.A(_009_),
    .Y(net91));
 BUFx2_ASAP7_75t_R rebuffer39 (.A(net91),
    .Y(net92));
 BUFx3_ASAP7_75t_R rebuffer40 (.A(_011_),
    .Y(net93));
 BUFx2_ASAP7_75t_R rebuffer41 (.A(net93),
    .Y(net94));
 BUFx2_ASAP7_75t_R rebuffer42 (.A(net94),
    .Y(net95));
 BUFx2_ASAP7_75t_R rebuffer43 (.A(net93),
    .Y(net96));
 BUFx2_ASAP7_75t_R rebuffer44 (.A(_101_),
    .Y(net97));
 BUFx2_ASAP7_75t_R rebuffer45 (.A(_291_),
    .Y(net98));
 BUFx2_ASAP7_75t_R rebuffer46 (.A(net98),
    .Y(net99));
 BUFx2_ASAP7_75t_R rebuffer47 (.A(\dpath.a_lt_b$in0[2] ),
    .Y(net100));
 BUFx2_ASAP7_75t_R rebuffer48 (.A(_030_),
    .Y(net101));
 BUFx3_ASAP7_75t_R rebuffer49 (.A(_097_),
    .Y(net102));
 BUFx2_ASAP7_75t_R rebuffer50 (.A(_296_),
    .Y(net103));
 BUFx2_ASAP7_75t_R rebuffer51 (.A(_007_),
    .Y(net104));
 BUFx3_ASAP7_75t_R rebuffer52 (.A(_007_),
    .Y(net105));
 BUFx2_ASAP7_75t_R rebuffer53 (.A(net105),
    .Y(net106));
 BUFx2_ASAP7_75t_R rebuffer36 (.A(_016_),
    .Y(net89));
 BUFx2_ASAP7_75t_R rebuffer54 (.A(_049_),
    .Y(net107));
 BUFx2_ASAP7_75t_R rebuffer58 (.A(_293_),
    .Y(net111));
 BUFx2_ASAP7_75t_R rebuffer59 (.A(_006_),
    .Y(net112));
 BUFx2_ASAP7_75t_R rebuffer60 (.A(_008_),
    .Y(net113));
 BUFx3_ASAP7_75t_R rebuffer61 (.A(net113),
    .Y(net114));
 OAI21x1_ASAP7_75t_R clone62 (.A1(_109_),
    .A2(_135_),
    .B(_136_),
    .Y(net115));
 BUFx2_ASAP7_75t_R clone63 (.A(_137_),
    .Y(net116));
 BUFx2_ASAP7_75t_R rebuffer64 (.A(_111_),
    .Y(net117));
 BUFx2_ASAP7_75t_R clone65 (.A(_137_),
    .Y(net118));
 BUFx2_ASAP7_75t_R clone66 (.A(_137_),
    .Y(net119));
 BUFx6f_ASAP7_75t_R rebuffer67 (.A(_137_),
    .Y(net120));
 BUFx2_ASAP7_75t_R rebuffer68 (.A(\dpath.a_lt_b$in0[8] ),
    .Y(net121));
 BUFx2_ASAP7_75t_R rebuffer69 (.A(_134_),
    .Y(net122));
 DECAPx10_ASAP7_75t_R FILLER_0_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46 ();
 DECAPx1_ASAP7_75t_R FILLER_0_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72 ();
 DECAPx6_ASAP7_75t_R FILLER_0_88 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144 ();
 FILLER_ASAP7_75t_R FILLER_0_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_174 ();
 DECAPx10_ASAP7_75t_R FILLER_0_196 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218 ();
 DECAPx6_ASAP7_75t_R FILLER_0_240 ();
 DECAPx1_ASAP7_75t_R FILLER_0_254 ();
 DECAPx10_ASAP7_75t_R FILLER_1_2 ();
 DECAPx10_ASAP7_75t_R FILLER_1_24 ();
 DECAPx10_ASAP7_75t_R FILLER_1_46 ();
 DECAPx10_ASAP7_75t_R FILLER_1_68 ();
 DECAPx10_ASAP7_75t_R FILLER_1_90 ();
 DECAPx10_ASAP7_75t_R FILLER_1_112 ();
 DECAPx10_ASAP7_75t_R FILLER_1_134 ();
 DECAPx10_ASAP7_75t_R FILLER_1_156 ();
 DECAPx10_ASAP7_75t_R FILLER_1_178 ();
 DECAPx10_ASAP7_75t_R FILLER_1_200 ();
 DECAPx10_ASAP7_75t_R FILLER_1_222 ();
 DECAPx6_ASAP7_75t_R FILLER_1_244 ();
 DECAPx10_ASAP7_75t_R FILLER_2_2 ();
 DECAPx10_ASAP7_75t_R FILLER_2_24 ();
 DECAPx10_ASAP7_75t_R FILLER_2_46 ();
 DECAPx10_ASAP7_75t_R FILLER_2_68 ();
 DECAPx10_ASAP7_75t_R FILLER_2_90 ();
 DECAPx10_ASAP7_75t_R FILLER_2_112 ();
 DECAPx10_ASAP7_75t_R FILLER_2_134 ();
 DECAPx10_ASAP7_75t_R FILLER_2_156 ();
 DECAPx10_ASAP7_75t_R FILLER_2_178 ();
 DECAPx10_ASAP7_75t_R FILLER_2_200 ();
 DECAPx10_ASAP7_75t_R FILLER_2_222 ();
 DECAPx6_ASAP7_75t_R FILLER_2_244 ();
 DECAPx10_ASAP7_75t_R FILLER_3_2 ();
 DECAPx10_ASAP7_75t_R FILLER_3_24 ();
 DECAPx10_ASAP7_75t_R FILLER_3_46 ();
 DECAPx10_ASAP7_75t_R FILLER_3_68 ();
 DECAPx10_ASAP7_75t_R FILLER_3_90 ();
 DECAPx10_ASAP7_75t_R FILLER_3_112 ();
 DECAPx10_ASAP7_75t_R FILLER_3_134 ();
 DECAPx10_ASAP7_75t_R FILLER_3_156 ();
 DECAPx10_ASAP7_75t_R FILLER_3_178 ();
 DECAPx10_ASAP7_75t_R FILLER_3_200 ();
 DECAPx10_ASAP7_75t_R FILLER_3_222 ();
 DECAPx6_ASAP7_75t_R FILLER_3_244 ();
 DECAPx10_ASAP7_75t_R FILLER_4_2 ();
 DECAPx10_ASAP7_75t_R FILLER_4_24 ();
 DECAPx10_ASAP7_75t_R FILLER_4_46 ();
 DECAPx10_ASAP7_75t_R FILLER_4_68 ();
 DECAPx10_ASAP7_75t_R FILLER_4_90 ();
 DECAPx10_ASAP7_75t_R FILLER_4_112 ();
 DECAPx10_ASAP7_75t_R FILLER_4_134 ();
 DECAPx10_ASAP7_75t_R FILLER_4_156 ();
 DECAPx10_ASAP7_75t_R FILLER_4_178 ();
 DECAPx10_ASAP7_75t_R FILLER_4_200 ();
 DECAPx10_ASAP7_75t_R FILLER_4_222 ();
 DECAPx6_ASAP7_75t_R FILLER_4_244 ();
 DECAPx10_ASAP7_75t_R FILLER_5_2 ();
 DECAPx10_ASAP7_75t_R FILLER_5_24 ();
 DECAPx10_ASAP7_75t_R FILLER_5_46 ();
 DECAPx10_ASAP7_75t_R FILLER_5_68 ();
 DECAPx10_ASAP7_75t_R FILLER_5_90 ();
 DECAPx10_ASAP7_75t_R FILLER_5_112 ();
 DECAPx10_ASAP7_75t_R FILLER_5_134 ();
 DECAPx10_ASAP7_75t_R FILLER_5_156 ();
 DECAPx10_ASAP7_75t_R FILLER_5_178 ();
 DECAPx10_ASAP7_75t_R FILLER_5_200 ();
 DECAPx10_ASAP7_75t_R FILLER_5_222 ();
 DECAPx6_ASAP7_75t_R FILLER_5_244 ();
 DECAPx10_ASAP7_75t_R FILLER_6_2 ();
 DECAPx10_ASAP7_75t_R FILLER_6_24 ();
 DECAPx10_ASAP7_75t_R FILLER_6_46 ();
 DECAPx10_ASAP7_75t_R FILLER_6_68 ();
 DECAPx10_ASAP7_75t_R FILLER_6_90 ();
 DECAPx10_ASAP7_75t_R FILLER_6_112 ();
 DECAPx10_ASAP7_75t_R FILLER_6_134 ();
 DECAPx10_ASAP7_75t_R FILLER_6_156 ();
 DECAPx10_ASAP7_75t_R FILLER_6_178 ();
 DECAPx10_ASAP7_75t_R FILLER_6_200 ();
 DECAPx10_ASAP7_75t_R FILLER_6_222 ();
 DECAPx6_ASAP7_75t_R FILLER_6_244 ();
 DECAPx10_ASAP7_75t_R FILLER_7_2 ();
 DECAPx10_ASAP7_75t_R FILLER_7_24 ();
 DECAPx10_ASAP7_75t_R FILLER_7_46 ();
 DECAPx10_ASAP7_75t_R FILLER_7_68 ();
 DECAPx10_ASAP7_75t_R FILLER_7_90 ();
 DECAPx10_ASAP7_75t_R FILLER_7_112 ();
 DECAPx10_ASAP7_75t_R FILLER_7_134 ();
 DECAPx10_ASAP7_75t_R FILLER_7_156 ();
 DECAPx10_ASAP7_75t_R FILLER_7_178 ();
 DECAPx10_ASAP7_75t_R FILLER_7_200 ();
 DECAPx10_ASAP7_75t_R FILLER_7_222 ();
 DECAPx6_ASAP7_75t_R FILLER_7_244 ();
 DECAPx10_ASAP7_75t_R FILLER_8_2 ();
 DECAPx10_ASAP7_75t_R FILLER_8_24 ();
 DECAPx10_ASAP7_75t_R FILLER_8_46 ();
 DECAPx10_ASAP7_75t_R FILLER_8_68 ();
 DECAPx10_ASAP7_75t_R FILLER_8_90 ();
 DECAPx10_ASAP7_75t_R FILLER_8_112 ();
 DECAPx10_ASAP7_75t_R FILLER_8_134 ();
 DECAPx10_ASAP7_75t_R FILLER_8_156 ();
 DECAPx10_ASAP7_75t_R FILLER_8_178 ();
 DECAPx10_ASAP7_75t_R FILLER_8_200 ();
 DECAPx10_ASAP7_75t_R FILLER_8_222 ();
 DECAPx6_ASAP7_75t_R FILLER_8_244 ();
 DECAPx10_ASAP7_75t_R FILLER_9_2 ();
 DECAPx10_ASAP7_75t_R FILLER_9_24 ();
 DECAPx10_ASAP7_75t_R FILLER_9_46 ();
 DECAPx10_ASAP7_75t_R FILLER_9_68 ();
 DECAPx10_ASAP7_75t_R FILLER_9_90 ();
 DECAPx10_ASAP7_75t_R FILLER_9_112 ();
 DECAPx10_ASAP7_75t_R FILLER_9_134 ();
 DECAPx10_ASAP7_75t_R FILLER_9_156 ();
 DECAPx10_ASAP7_75t_R FILLER_9_178 ();
 DECAPx10_ASAP7_75t_R FILLER_9_200 ();
 DECAPx10_ASAP7_75t_R FILLER_9_222 ();
 DECAPx6_ASAP7_75t_R FILLER_9_244 ();
 DECAPx10_ASAP7_75t_R FILLER_10_2 ();
 DECAPx10_ASAP7_75t_R FILLER_10_24 ();
 DECAPx10_ASAP7_75t_R FILLER_10_46 ();
 DECAPx10_ASAP7_75t_R FILLER_10_68 ();
 DECAPx10_ASAP7_75t_R FILLER_10_90 ();
 DECAPx10_ASAP7_75t_R FILLER_10_112 ();
 DECAPx10_ASAP7_75t_R FILLER_10_134 ();
 DECAPx10_ASAP7_75t_R FILLER_10_156 ();
 DECAPx10_ASAP7_75t_R FILLER_10_178 ();
 DECAPx10_ASAP7_75t_R FILLER_10_200 ();
 DECAPx10_ASAP7_75t_R FILLER_10_222 ();
 DECAPx6_ASAP7_75t_R FILLER_10_244 ();
 DECAPx6_ASAP7_75t_R FILLER_11_2 ();
 DECAPx10_ASAP7_75t_R FILLER_11_21 ();
 DECAPx10_ASAP7_75t_R FILLER_11_43 ();
 DECAPx4_ASAP7_75t_R FILLER_11_65 ();
 FILLER_ASAP7_75t_R FILLER_11_75 ();
 DECAPx10_ASAP7_75t_R FILLER_11_83 ();
 DECAPx10_ASAP7_75t_R FILLER_11_105 ();
 DECAPx10_ASAP7_75t_R FILLER_11_127 ();
 DECAPx10_ASAP7_75t_R FILLER_11_149 ();
 DECAPx10_ASAP7_75t_R FILLER_11_171 ();
 DECAPx10_ASAP7_75t_R FILLER_11_193 ();
 DECAPx10_ASAP7_75t_R FILLER_11_215 ();
 DECAPx6_ASAP7_75t_R FILLER_11_237 ();
 DECAPx2_ASAP7_75t_R FILLER_11_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_257 ();
 DECAPx10_ASAP7_75t_R FILLER_12_2 ();
 DECAPx4_ASAP7_75t_R FILLER_12_24 ();
 FILLER_ASAP7_75t_R FILLER_12_34 ();
 DECAPx10_ASAP7_75t_R FILLER_12_42 ();
 DECAPx2_ASAP7_75t_R FILLER_12_64 ();
 FILLER_ASAP7_75t_R FILLER_12_70 ();
 FILLER_ASAP7_75t_R FILLER_12_93 ();
 DECAPx6_ASAP7_75t_R FILLER_12_101 ();
 DECAPx10_ASAP7_75t_R FILLER_12_142 ();
 DECAPx10_ASAP7_75t_R FILLER_12_164 ();
 DECAPx10_ASAP7_75t_R FILLER_12_186 ();
 DECAPx10_ASAP7_75t_R FILLER_12_208 ();
 DECAPx10_ASAP7_75t_R FILLER_12_230 ();
 DECAPx2_ASAP7_75t_R FILLER_12_252 ();
 DECAPx10_ASAP7_75t_R FILLER_13_2 ();
 DECAPx10_ASAP7_75t_R FILLER_13_24 ();
 FILLER_ASAP7_75t_R FILLER_13_75 ();
 DECAPx6_ASAP7_75t_R FILLER_13_85 ();
 DECAPx6_ASAP7_75t_R FILLER_13_128 ();
 DECAPx10_ASAP7_75t_R FILLER_13_163 ();
 DECAPx10_ASAP7_75t_R FILLER_13_185 ();
 DECAPx10_ASAP7_75t_R FILLER_13_207 ();
 DECAPx10_ASAP7_75t_R FILLER_13_229 ();
 DECAPx2_ASAP7_75t_R FILLER_13_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_257 ();
 DECAPx10_ASAP7_75t_R FILLER_14_2 ();
 DECAPx1_ASAP7_75t_R FILLER_14_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_28 ();
 DECAPx6_ASAP7_75t_R FILLER_14_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_51 ();
 DECAPx6_ASAP7_75t_R FILLER_14_58 ();
 DECAPx1_ASAP7_75t_R FILLER_14_72 ();
 DECAPx4_ASAP7_75t_R FILLER_14_82 ();
 DECAPx6_ASAP7_75t_R FILLER_14_106 ();
 FILLER_ASAP7_75t_R FILLER_14_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_122 ();
 DECAPx6_ASAP7_75t_R FILLER_14_129 ();
 DECAPx1_ASAP7_75t_R FILLER_14_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_147 ();
 DECAPx10_ASAP7_75t_R FILLER_14_154 ();
 DECAPx10_ASAP7_75t_R FILLER_14_176 ();
 DECAPx10_ASAP7_75t_R FILLER_14_198 ();
 DECAPx10_ASAP7_75t_R FILLER_14_220 ();
 DECAPx6_ASAP7_75t_R FILLER_14_242 ();
 FILLER_ASAP7_75t_R FILLER_14_256 ();
 DECAPx10_ASAP7_75t_R FILLER_15_2 ();
 DECAPx6_ASAP7_75t_R FILLER_15_24 ();
 FILLER_ASAP7_75t_R FILLER_15_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_40 ();
 DECAPx1_ASAP7_75t_R FILLER_15_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_73 ();
 DECAPx6_ASAP7_75t_R FILLER_15_80 ();
 DECAPx2_ASAP7_75t_R FILLER_15_94 ();
 DECAPx10_ASAP7_75t_R FILLER_15_106 ();
 DECAPx6_ASAP7_75t_R FILLER_15_128 ();
 DECAPx2_ASAP7_75t_R FILLER_15_156 ();
 FILLER_ASAP7_75t_R FILLER_15_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_164 ();
 DECAPx10_ASAP7_75t_R FILLER_15_186 ();
 DECAPx10_ASAP7_75t_R FILLER_15_208 ();
 DECAPx10_ASAP7_75t_R FILLER_15_230 ();
 DECAPx2_ASAP7_75t_R FILLER_15_252 ();
 DECAPx10_ASAP7_75t_R FILLER_16_2 ();
 DECAPx2_ASAP7_75t_R FILLER_16_24 ();
 FILLER_ASAP7_75t_R FILLER_16_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_51 ();
 DECAPx6_ASAP7_75t_R FILLER_16_58 ();
 DECAPx2_ASAP7_75t_R FILLER_16_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_89 ();
 DECAPx4_ASAP7_75t_R FILLER_16_112 ();
 FILLER_ASAP7_75t_R FILLER_16_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_124 ();
 DECAPx6_ASAP7_75t_R FILLER_16_131 ();
 DECAPx2_ASAP7_75t_R FILLER_16_145 ();
 DECAPx10_ASAP7_75t_R FILLER_16_160 ();
 DECAPx10_ASAP7_75t_R FILLER_16_182 ();
 DECAPx2_ASAP7_75t_R FILLER_16_204 ();
 DECAPx10_ASAP7_75t_R FILLER_16_216 ();
 DECAPx6_ASAP7_75t_R FILLER_16_238 ();
 DECAPx2_ASAP7_75t_R FILLER_16_252 ();
 DECAPx6_ASAP7_75t_R FILLER_17_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_16 ();
 DECAPx10_ASAP7_75t_R FILLER_17_22 ();
 DECAPx10_ASAP7_75t_R FILLER_17_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_66 ();
 DECAPx6_ASAP7_75t_R FILLER_17_89 ();
 DECAPx1_ASAP7_75t_R FILLER_17_103 ();
 DECAPx4_ASAP7_75t_R FILLER_17_117 ();
 FILLER_ASAP7_75t_R FILLER_17_127 ();
 DECAPx10_ASAP7_75t_R FILLER_17_133 ();
 FILLER_ASAP7_75t_R FILLER_17_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_157 ();
 DECAPx4_ASAP7_75t_R FILLER_17_170 ();
 DECAPx1_ASAP7_75t_R FILLER_17_224 ();
 DECAPx10_ASAP7_75t_R FILLER_17_233 ();
 FILLER_ASAP7_75t_R FILLER_17_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_257 ();
 DECAPx10_ASAP7_75t_R FILLER_18_2 ();
 DECAPx6_ASAP7_75t_R FILLER_18_24 ();
 DECAPx2_ASAP7_75t_R FILLER_18_64 ();
 FILLER_ASAP7_75t_R FILLER_18_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_72 ();
 DECAPx1_ASAP7_75t_R FILLER_18_79 ();
 DECAPx6_ASAP7_75t_R FILLER_18_91 ();
 FILLER_ASAP7_75t_R FILLER_18_105 ();
 DECAPx1_ASAP7_75t_R FILLER_18_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_117 ();
 DECAPx2_ASAP7_75t_R FILLER_18_146 ();
 FILLER_ASAP7_75t_R FILLER_18_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_163 ();
 DECAPx6_ASAP7_75t_R FILLER_18_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_190 ();
 DECAPx10_ASAP7_75t_R FILLER_18_212 ();
 DECAPx10_ASAP7_75t_R FILLER_18_234 ();
 FILLER_ASAP7_75t_R FILLER_18_256 ();
 DECAPx10_ASAP7_75t_R FILLER_19_2 ();
 DECAPx10_ASAP7_75t_R FILLER_19_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_46 ();
 DECAPx2_ASAP7_75t_R FILLER_19_65 ();
 FILLER_ASAP7_75t_R FILLER_19_71 ();
 DECAPx2_ASAP7_75t_R FILLER_19_89 ();
 FILLER_ASAP7_75t_R FILLER_19_95 ();
 DECAPx4_ASAP7_75t_R FILLER_19_113 ();
 DECAPx6_ASAP7_75t_R FILLER_19_139 ();
 DECAPx2_ASAP7_75t_R FILLER_19_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_159 ();
 DECAPx10_ASAP7_75t_R FILLER_19_168 ();
 DECAPx2_ASAP7_75t_R FILLER_19_190 ();
 DECAPx10_ASAP7_75t_R FILLER_19_202 ();
 DECAPx10_ASAP7_75t_R FILLER_19_224 ();
 DECAPx4_ASAP7_75t_R FILLER_19_246 ();
 FILLER_ASAP7_75t_R FILLER_19_256 ();
 DECAPx10_ASAP7_75t_R FILLER_20_2 ();
 DECAPx6_ASAP7_75t_R FILLER_20_24 ();
 DECAPx2_ASAP7_75t_R FILLER_20_38 ();
 FILLER_ASAP7_75t_R FILLER_20_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_76 ();
 DECAPx10_ASAP7_75t_R FILLER_20_83 ();
 DECAPx6_ASAP7_75t_R FILLER_20_105 ();
 DECAPx2_ASAP7_75t_R FILLER_20_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_125 ();
 DECAPx10_ASAP7_75t_R FILLER_20_132 ();
 FILLER_ASAP7_75t_R FILLER_20_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_156 ();
 DECAPx6_ASAP7_75t_R FILLER_20_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_179 ();
 DECAPx2_ASAP7_75t_R FILLER_20_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_195 ();
 DECAPx1_ASAP7_75t_R FILLER_20_204 ();
 DECAPx10_ASAP7_75t_R FILLER_20_214 ();
 DECAPx10_ASAP7_75t_R FILLER_20_236 ();
 DECAPx1_ASAP7_75t_R FILLER_21_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_6 ();
 DECAPx1_ASAP7_75t_R FILLER_21_12 ();
 FILLER_ASAP7_75t_R FILLER_21_22 ();
 DECAPx10_ASAP7_75t_R FILLER_21_35 ();
 FILLER_ASAP7_75t_R FILLER_21_57 ();
 DECAPx2_ASAP7_75t_R FILLER_21_65 ();
 FILLER_ASAP7_75t_R FILLER_21_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_73 ();
 DECAPx6_ASAP7_75t_R FILLER_21_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_98 ();
 DECAPx6_ASAP7_75t_R FILLER_21_105 ();
 DECAPx1_ASAP7_75t_R FILLER_21_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_123 ();
 DECAPx4_ASAP7_75t_R FILLER_21_133 ();
 FILLER_ASAP7_75t_R FILLER_21_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_145 ();
 DECAPx1_ASAP7_75t_R FILLER_21_153 ();
 DECAPx1_ASAP7_75t_R FILLER_21_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_167 ();
 DECAPx2_ASAP7_75t_R FILLER_21_174 ();
 FILLER_ASAP7_75t_R FILLER_21_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_182 ();
 FILLER_ASAP7_75t_R FILLER_21_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_197 ();
 DECAPx10_ASAP7_75t_R FILLER_21_206 ();
 DECAPx10_ASAP7_75t_R FILLER_21_228 ();
 DECAPx2_ASAP7_75t_R FILLER_21_250 ();
 FILLER_ASAP7_75t_R FILLER_21_256 ();
 DECAPx1_ASAP7_75t_R FILLER_22_2 ();
 DECAPx6_ASAP7_75t_R FILLER_22_11 ();
 DECAPx1_ASAP7_75t_R FILLER_22_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_29 ();
 DECAPx6_ASAP7_75t_R FILLER_22_44 ();
 DECAPx2_ASAP7_75t_R FILLER_22_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_64 ();
 DECAPx1_ASAP7_75t_R FILLER_22_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_92 ();
 DECAPx2_ASAP7_75t_R FILLER_22_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_116 ();
 FILLER_ASAP7_75t_R FILLER_22_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_131 ();
 DECAPx4_ASAP7_75t_R FILLER_22_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_148 ();
 DECAPx1_ASAP7_75t_R FILLER_22_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_171 ();
 DECAPx6_ASAP7_75t_R FILLER_22_178 ();
 FILLER_ASAP7_75t_R FILLER_22_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_194 ();
 DECAPx2_ASAP7_75t_R FILLER_22_200 ();
 FILLER_ASAP7_75t_R FILLER_22_206 ();
 DECAPx6_ASAP7_75t_R FILLER_22_222 ();
 DECAPx1_ASAP7_75t_R FILLER_22_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_240 ();
 DECAPx4_ASAP7_75t_R FILLER_22_246 ();
 FILLER_ASAP7_75t_R FILLER_22_256 ();
 DECAPx4_ASAP7_75t_R FILLER_23_2 ();
 DECAPx2_ASAP7_75t_R FILLER_23_33 ();
 DECAPx4_ASAP7_75t_R FILLER_23_51 ();
 FILLER_ASAP7_75t_R FILLER_23_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_63 ();
 FILLER_ASAP7_75t_R FILLER_23_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_78 ();
 FILLER_ASAP7_75t_R FILLER_23_91 ();
 DECAPx10_ASAP7_75t_R FILLER_23_119 ();
 DECAPx2_ASAP7_75t_R FILLER_23_141 ();
 FILLER_ASAP7_75t_R FILLER_23_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_149 ();
 DECAPx2_ASAP7_75t_R FILLER_23_172 ();
 FILLER_ASAP7_75t_R FILLER_23_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_180 ();
 DECAPx6_ASAP7_75t_R FILLER_23_222 ();
 DECAPx1_ASAP7_75t_R FILLER_23_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_240 ();
 FILLER_ASAP7_75t_R FILLER_23_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_248 ();
 DECAPx1_ASAP7_75t_R FILLER_23_254 ();
 DECAPx6_ASAP7_75t_R FILLER_24_2 ();
 DECAPx1_ASAP7_75t_R FILLER_24_16 ();
 DECAPx4_ASAP7_75t_R FILLER_24_25 ();
 FILLER_ASAP7_75t_R FILLER_24_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_53 ();
 FILLER_ASAP7_75t_R FILLER_24_60 ();
 FILLER_ASAP7_75t_R FILLER_24_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_79 ();
 DECAPx6_ASAP7_75t_R FILLER_24_127 ();
 DECAPx1_ASAP7_75t_R FILLER_24_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_153 ();
 DECAPx1_ASAP7_75t_R FILLER_24_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_166 ();
 DECAPx2_ASAP7_75t_R FILLER_24_174 ();
 FILLER_ASAP7_75t_R FILLER_24_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_182 ();
 DECAPx4_ASAP7_75t_R FILLER_24_199 ();
 FILLER_ASAP7_75t_R FILLER_24_209 ();
 DECAPx10_ASAP7_75t_R FILLER_24_217 ();
 DECAPx6_ASAP7_75t_R FILLER_24_239 ();
 DECAPx1_ASAP7_75t_R FILLER_24_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_257 ();
 DECAPx10_ASAP7_75t_R FILLER_25_2 ();
 DECAPx1_ASAP7_75t_R FILLER_25_24 ();
 DECAPx6_ASAP7_75t_R FILLER_25_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_92 ();
 DECAPx6_ASAP7_75t_R FILLER_25_127 ();
 DECAPx2_ASAP7_75t_R FILLER_25_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_182 ();
 DECAPx1_ASAP7_75t_R FILLER_25_194 ();
 DECAPx10_ASAP7_75t_R FILLER_25_212 ();
 DECAPx10_ASAP7_75t_R FILLER_25_234 ();
 FILLER_ASAP7_75t_R FILLER_25_256 ();
 DECAPx6_ASAP7_75t_R FILLER_26_2 ();
 FILLER_ASAP7_75t_R FILLER_26_16 ();
 DECAPx6_ASAP7_75t_R FILLER_26_23 ();
 DECAPx2_ASAP7_75t_R FILLER_26_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_43 ();
 DECAPx1_ASAP7_75t_R FILLER_26_53 ();
 FILLER_ASAP7_75t_R FILLER_26_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_89 ();
 DECAPx6_ASAP7_75t_R FILLER_26_96 ();
 FILLER_ASAP7_75t_R FILLER_26_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_112 ();
 DECAPx10_ASAP7_75t_R FILLER_26_129 ();
 DECAPx2_ASAP7_75t_R FILLER_26_151 ();
 FILLER_ASAP7_75t_R FILLER_26_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_185 ();
 DECAPx2_ASAP7_75t_R FILLER_26_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_204 ();
 DECAPx10_ASAP7_75t_R FILLER_26_226 ();
 DECAPx4_ASAP7_75t_R FILLER_26_248 ();
 DECAPx10_ASAP7_75t_R FILLER_27_2 ();
 DECAPx4_ASAP7_75t_R FILLER_27_24 ();
 FILLER_ASAP7_75t_R FILLER_27_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_36 ();
 DECAPx1_ASAP7_75t_R FILLER_27_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_47 ();
 FILLER_ASAP7_75t_R FILLER_27_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_61 ();
 FILLER_ASAP7_75t_R FILLER_27_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_70 ();
 DECAPx6_ASAP7_75t_R FILLER_27_100 ();
 DECAPx1_ASAP7_75t_R FILLER_27_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_125 ();
 FILLER_ASAP7_75t_R FILLER_27_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_140 ();
 FILLER_ASAP7_75t_R FILLER_27_144 ();
 DECAPx1_ASAP7_75t_R FILLER_27_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_157 ();
 DECAPx1_ASAP7_75t_R FILLER_27_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_199 ();
 DECAPx6_ASAP7_75t_R FILLER_27_214 ();
 FILLER_ASAP7_75t_R FILLER_27_228 ();
 DECAPx10_ASAP7_75t_R FILLER_27_236 ();
 FILLER_ASAP7_75t_R FILLER_28_2 ();
 DECAPx4_ASAP7_75t_R FILLER_28_14 ();
 FILLER_ASAP7_75t_R FILLER_28_24 ();
 DECAPx10_ASAP7_75t_R FILLER_28_53 ();
 DECAPx10_ASAP7_75t_R FILLER_28_80 ();
 DECAPx6_ASAP7_75t_R FILLER_28_102 ();
 DECAPx1_ASAP7_75t_R FILLER_28_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_128 ();
 DECAPx2_ASAP7_75t_R FILLER_28_162 ();
 FILLER_ASAP7_75t_R FILLER_28_168 ();
 FILLER_ASAP7_75t_R FILLER_28_173 ();
 DECAPx1_ASAP7_75t_R FILLER_28_189 ();
 DECAPx10_ASAP7_75t_R FILLER_28_205 ();
 DECAPx1_ASAP7_75t_R FILLER_28_227 ();
 DECAPx10_ASAP7_75t_R FILLER_28_236 ();
 DECAPx1_ASAP7_75t_R FILLER_29_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_6 ();
 DECAPx2_ASAP7_75t_R FILLER_29_28 ();
 FILLER_ASAP7_75t_R FILLER_29_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_60 ();
 DECAPx10_ASAP7_75t_R FILLER_29_68 ();
 DECAPx10_ASAP7_75t_R FILLER_29_90 ();
 FILLER_ASAP7_75t_R FILLER_29_117 ();
 DECAPx1_ASAP7_75t_R FILLER_29_131 ();
 FILLER_ASAP7_75t_R FILLER_29_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_148 ();
 FILLER_ASAP7_75t_R FILLER_29_162 ();
 FILLER_ASAP7_75t_R FILLER_29_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_182 ();
 DECAPx10_ASAP7_75t_R FILLER_29_200 ();
 DECAPx10_ASAP7_75t_R FILLER_29_222 ();
 DECAPx6_ASAP7_75t_R FILLER_29_244 ();
 DECAPx6_ASAP7_75t_R FILLER_30_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_62 ();
 FILLER_ASAP7_75t_R FILLER_30_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_77 ();
 DECAPx10_ASAP7_75t_R FILLER_30_83 ();
 DECAPx4_ASAP7_75t_R FILLER_30_105 ();
 DECAPx2_ASAP7_75t_R FILLER_30_121 ();
 DECAPx6_ASAP7_75t_R FILLER_30_136 ();
 FILLER_ASAP7_75t_R FILLER_30_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_157 ();
 FILLER_ASAP7_75t_R FILLER_30_163 ();
 DECAPx6_ASAP7_75t_R FILLER_30_176 ();
 DECAPx1_ASAP7_75t_R FILLER_30_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_194 ();
 DECAPx6_ASAP7_75t_R FILLER_30_207 ();
 DECAPx2_ASAP7_75t_R FILLER_30_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_227 ();
 DECAPx10_ASAP7_75t_R FILLER_30_233 ();
 FILLER_ASAP7_75t_R FILLER_30_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_257 ();
 DECAPx10_ASAP7_75t_R FILLER_31_2 ();
 DECAPx2_ASAP7_75t_R FILLER_31_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_30 ();
 FILLER_ASAP7_75t_R FILLER_31_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_41 ();
 DECAPx6_ASAP7_75t_R FILLER_31_71 ();
 DECAPx2_ASAP7_75t_R FILLER_31_85 ();
 DECAPx10_ASAP7_75t_R FILLER_31_101 ();
 DECAPx10_ASAP7_75t_R FILLER_31_123 ();
 DECAPx10_ASAP7_75t_R FILLER_31_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_167 ();
 DECAPx10_ASAP7_75t_R FILLER_31_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_196 ();
 DECAPx10_ASAP7_75t_R FILLER_31_208 ();
 DECAPx10_ASAP7_75t_R FILLER_31_230 ();
 DECAPx2_ASAP7_75t_R FILLER_31_252 ();
 DECAPx4_ASAP7_75t_R FILLER_32_2 ();
 DECAPx6_ASAP7_75t_R FILLER_32_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_42 ();
 FILLER_ASAP7_75t_R FILLER_32_66 ();
 DECAPx4_ASAP7_75t_R FILLER_32_76 ();
 FILLER_ASAP7_75t_R FILLER_32_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_88 ();
 DECAPx6_ASAP7_75t_R FILLER_32_102 ();
 DECAPx1_ASAP7_75t_R FILLER_32_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_120 ();
 DECAPx10_ASAP7_75t_R FILLER_32_131 ();
 DECAPx6_ASAP7_75t_R FILLER_32_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_167 ();
 DECAPx2_ASAP7_75t_R FILLER_32_183 ();
 DECAPx4_ASAP7_75t_R FILLER_32_198 ();
 FILLER_ASAP7_75t_R FILLER_32_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_217 ();
 DECAPx2_ASAP7_75t_R FILLER_32_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_230 ();
 DECAPx10_ASAP7_75t_R FILLER_32_236 ();
 FILLER_ASAP7_75t_R FILLER_33_2 ();
 DECAPx6_ASAP7_75t_R FILLER_33_9 ();
 FILLER_ASAP7_75t_R FILLER_33_23 ();
 DECAPx4_ASAP7_75t_R FILLER_33_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_41 ();
 FILLER_ASAP7_75t_R FILLER_33_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_51 ();
 FILLER_ASAP7_75t_R FILLER_33_62 ();
 DECAPx2_ASAP7_75t_R FILLER_33_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_83 ();
 FILLER_ASAP7_75t_R FILLER_33_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_123 ();
 DECAPx10_ASAP7_75t_R FILLER_33_127 ();
 DECAPx4_ASAP7_75t_R FILLER_33_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_159 ();
 DECAPx2_ASAP7_75t_R FILLER_33_174 ();
 FILLER_ASAP7_75t_R FILLER_33_180 ();
 DECAPx6_ASAP7_75t_R FILLER_33_188 ();
 DECAPx2_ASAP7_75t_R FILLER_33_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_208 ();
 DECAPx6_ASAP7_75t_R FILLER_33_238 ();
 DECAPx2_ASAP7_75t_R FILLER_33_252 ();
 DECAPx1_ASAP7_75t_R FILLER_34_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_6 ();
 FILLER_ASAP7_75t_R FILLER_34_12 ();
 DECAPx2_ASAP7_75t_R FILLER_34_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_41 ();
 DECAPx2_ASAP7_75t_R FILLER_34_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_57 ();
 DECAPx10_ASAP7_75t_R FILLER_34_70 ();
 DECAPx1_ASAP7_75t_R FILLER_34_92 ();
 FILLER_ASAP7_75t_R FILLER_34_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_104 ();
 DECAPx2_ASAP7_75t_R FILLER_34_133 ();
 DECAPx10_ASAP7_75t_R FILLER_34_153 ();
 DECAPx10_ASAP7_75t_R FILLER_34_175 ();
 FILLER_ASAP7_75t_R FILLER_34_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_207 ();
 DECAPx1_ASAP7_75t_R FILLER_34_211 ();
 DECAPx2_ASAP7_75t_R FILLER_34_221 ();
 FILLER_ASAP7_75t_R FILLER_34_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_229 ();
 DECAPx10_ASAP7_75t_R FILLER_34_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_257 ();
 DECAPx10_ASAP7_75t_R FILLER_35_2 ();
 FILLER_ASAP7_75t_R FILLER_35_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_26 ();
 FILLER_ASAP7_75t_R FILLER_35_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_37 ();
 FILLER_ASAP7_75t_R FILLER_35_56 ();
 DECAPx4_ASAP7_75t_R FILLER_35_73 ();
 FILLER_ASAP7_75t_R FILLER_35_83 ();
 DECAPx10_ASAP7_75t_R FILLER_35_93 ();
 DECAPx1_ASAP7_75t_R FILLER_35_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_119 ();
 DECAPx6_ASAP7_75t_R FILLER_35_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_158 ();
 DECAPx6_ASAP7_75t_R FILLER_35_180 ();
 DECAPx2_ASAP7_75t_R FILLER_35_194 ();
 FILLER_ASAP7_75t_R FILLER_35_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_216 ();
 DECAPx1_ASAP7_75t_R FILLER_35_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_227 ();
 DECAPx10_ASAP7_75t_R FILLER_35_233 ();
 FILLER_ASAP7_75t_R FILLER_35_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_257 ();
 FILLER_ASAP7_75t_R FILLER_36_2 ();
 DECAPx1_ASAP7_75t_R FILLER_36_47 ();
 DECAPx10_ASAP7_75t_R FILLER_36_66 ();
 DECAPx10_ASAP7_75t_R FILLER_36_88 ();
 DECAPx4_ASAP7_75t_R FILLER_36_110 ();
 FILLER_ASAP7_75t_R FILLER_36_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_122 ();
 DECAPx6_ASAP7_75t_R FILLER_36_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_164 ();
 DECAPx6_ASAP7_75t_R FILLER_36_178 ();
 DECAPx1_ASAP7_75t_R FILLER_36_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_196 ();
 DECAPx10_ASAP7_75t_R FILLER_36_218 ();
 DECAPx6_ASAP7_75t_R FILLER_36_240 ();
 DECAPx1_ASAP7_75t_R FILLER_36_254 ();
 DECAPx6_ASAP7_75t_R FILLER_37_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_16 ();
 DECAPx2_ASAP7_75t_R FILLER_37_27 ();
 DECAPx4_ASAP7_75t_R FILLER_37_39 ();
 DECAPx10_ASAP7_75t_R FILLER_37_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_99 ();
 DECAPx10_ASAP7_75t_R FILLER_37_120 ();
 DECAPx6_ASAP7_75t_R FILLER_37_142 ();
 DECAPx2_ASAP7_75t_R FILLER_37_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_170 ();
 DECAPx10_ASAP7_75t_R FILLER_37_183 ();
 DECAPx10_ASAP7_75t_R FILLER_37_205 ();
 DECAPx10_ASAP7_75t_R FILLER_37_227 ();
 DECAPx2_ASAP7_75t_R FILLER_37_249 ();
 FILLER_ASAP7_75t_R FILLER_37_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_257 ();
 DECAPx10_ASAP7_75t_R FILLER_38_2 ();
 DECAPx10_ASAP7_75t_R FILLER_38_24 ();
 DECAPx4_ASAP7_75t_R FILLER_38_46 ();
 FILLER_ASAP7_75t_R FILLER_38_56 ();
 DECAPx6_ASAP7_75t_R FILLER_38_64 ();
 DECAPx1_ASAP7_75t_R FILLER_38_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_82 ();
 DECAPx10_ASAP7_75t_R FILLER_38_91 ();
 DECAPx1_ASAP7_75t_R FILLER_38_113 ();
 DECAPx4_ASAP7_75t_R FILLER_38_125 ();
 FILLER_ASAP7_75t_R FILLER_38_135 ();
 DECAPx1_ASAP7_75t_R FILLER_38_145 ();
 DECAPx6_ASAP7_75t_R FILLER_38_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_179 ();
 DECAPx10_ASAP7_75t_R FILLER_38_200 ();
 DECAPx10_ASAP7_75t_R FILLER_38_222 ();
 DECAPx6_ASAP7_75t_R FILLER_38_244 ();
 DECAPx10_ASAP7_75t_R FILLER_39_2 ();
 DECAPx10_ASAP7_75t_R FILLER_39_24 ();
 DECAPx1_ASAP7_75t_R FILLER_39_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_50 ();
 DECAPx2_ASAP7_75t_R FILLER_39_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_65 ();
 FILLER_ASAP7_75t_R FILLER_39_72 ();
 DECAPx10_ASAP7_75t_R FILLER_39_80 ();
 DECAPx10_ASAP7_75t_R FILLER_39_102 ();
 DECAPx10_ASAP7_75t_R FILLER_39_124 ();
 FILLER_ASAP7_75t_R FILLER_39_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_148 ();
 DECAPx6_ASAP7_75t_R FILLER_39_155 ();
 DECAPx2_ASAP7_75t_R FILLER_39_169 ();
 DECAPx10_ASAP7_75t_R FILLER_39_196 ();
 DECAPx10_ASAP7_75t_R FILLER_39_218 ();
 DECAPx6_ASAP7_75t_R FILLER_39_240 ();
 DECAPx1_ASAP7_75t_R FILLER_39_254 ();
 DECAPx10_ASAP7_75t_R FILLER_40_2 ();
 DECAPx6_ASAP7_75t_R FILLER_40_24 ();
 DECAPx1_ASAP7_75t_R FILLER_40_38 ();
 DECAPx10_ASAP7_75t_R FILLER_40_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_70 ();
 DECAPx10_ASAP7_75t_R FILLER_40_87 ();
 FILLER_ASAP7_75t_R FILLER_40_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_111 ();
 DECAPx6_ASAP7_75t_R FILLER_40_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_151 ();
 DECAPx10_ASAP7_75t_R FILLER_40_158 ();
 DECAPx10_ASAP7_75t_R FILLER_40_180 ();
 DECAPx10_ASAP7_75t_R FILLER_40_202 ();
 DECAPx10_ASAP7_75t_R FILLER_40_224 ();
 DECAPx4_ASAP7_75t_R FILLER_40_246 ();
 FILLER_ASAP7_75t_R FILLER_40_256 ();
 DECAPx10_ASAP7_75t_R FILLER_41_2 ();
 DECAPx6_ASAP7_75t_R FILLER_41_24 ();
 FILLER_ASAP7_75t_R FILLER_41_38 ();
 DECAPx4_ASAP7_75t_R FILLER_41_50 ();
 FILLER_ASAP7_75t_R FILLER_41_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_62 ();
 FILLER_ASAP7_75t_R FILLER_41_89 ();
 DECAPx6_ASAP7_75t_R FILLER_41_97 ();
 DECAPx2_ASAP7_75t_R FILLER_41_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_117 ();
 DECAPx2_ASAP7_75t_R FILLER_41_134 ();
 DECAPx6_ASAP7_75t_R FILLER_41_177 ();
 DECAPx2_ASAP7_75t_R FILLER_41_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_197 ();
 DECAPx10_ASAP7_75t_R FILLER_41_206 ();
 DECAPx10_ASAP7_75t_R FILLER_41_228 ();
 DECAPx2_ASAP7_75t_R FILLER_41_250 ();
 FILLER_ASAP7_75t_R FILLER_41_256 ();
 DECAPx6_ASAP7_75t_R FILLER_42_2 ();
 FILLER_ASAP7_75t_R FILLER_42_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_18 ();
 FILLER_ASAP7_75t_R FILLER_42_40 ();
 FILLER_ASAP7_75t_R FILLER_42_65 ();
 DECAPx4_ASAP7_75t_R FILLER_42_87 ();
 DECAPx1_ASAP7_75t_R FILLER_42_103 ();
 DECAPx6_ASAP7_75t_R FILLER_42_134 ();
 DECAPx1_ASAP7_75t_R FILLER_42_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_159 ();
 DECAPx10_ASAP7_75t_R FILLER_42_200 ();
 DECAPx10_ASAP7_75t_R FILLER_42_222 ();
 DECAPx6_ASAP7_75t_R FILLER_42_244 ();
 DECAPx10_ASAP7_75t_R FILLER_43_2 ();
 DECAPx2_ASAP7_75t_R FILLER_43_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_30 ();
 DECAPx1_ASAP7_75t_R FILLER_43_58 ();
 DECAPx10_ASAP7_75t_R FILLER_43_95 ();
 DECAPx1_ASAP7_75t_R FILLER_43_117 ();
 FILLER_ASAP7_75t_R FILLER_43_161 ();
 FILLER_ASAP7_75t_R FILLER_43_166 ();
 DECAPx10_ASAP7_75t_R FILLER_43_189 ();
 DECAPx10_ASAP7_75t_R FILLER_43_211 ();
 DECAPx10_ASAP7_75t_R FILLER_43_233 ();
 FILLER_ASAP7_75t_R FILLER_43_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_257 ();
 DECAPx10_ASAP7_75t_R FILLER_44_2 ();
 DECAPx10_ASAP7_75t_R FILLER_44_24 ();
 DECAPx10_ASAP7_75t_R FILLER_44_46 ();
 DECAPx6_ASAP7_75t_R FILLER_44_68 ();
 FILLER_ASAP7_75t_R FILLER_44_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_84 ();
 DECAPx6_ASAP7_75t_R FILLER_44_106 ();
 DECAPx2_ASAP7_75t_R FILLER_44_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_126 ();
 DECAPx10_ASAP7_75t_R FILLER_44_154 ();
 DECAPx10_ASAP7_75t_R FILLER_44_176 ();
 DECAPx10_ASAP7_75t_R FILLER_44_198 ();
 DECAPx10_ASAP7_75t_R FILLER_44_220 ();
 DECAPx6_ASAP7_75t_R FILLER_44_242 ();
 FILLER_ASAP7_75t_R FILLER_44_256 ();
 DECAPx10_ASAP7_75t_R FILLER_45_2 ();
 DECAPx10_ASAP7_75t_R FILLER_45_24 ();
 DECAPx10_ASAP7_75t_R FILLER_45_46 ();
 DECAPx10_ASAP7_75t_R FILLER_45_68 ();
 DECAPx10_ASAP7_75t_R FILLER_45_90 ();
 DECAPx10_ASAP7_75t_R FILLER_45_112 ();
 DECAPx10_ASAP7_75t_R FILLER_45_134 ();
 DECAPx10_ASAP7_75t_R FILLER_45_156 ();
 DECAPx10_ASAP7_75t_R FILLER_45_178 ();
 DECAPx10_ASAP7_75t_R FILLER_45_200 ();
 DECAPx10_ASAP7_75t_R FILLER_45_222 ();
 DECAPx6_ASAP7_75t_R FILLER_45_244 ();
 DECAPx10_ASAP7_75t_R FILLER_46_2 ();
 DECAPx10_ASAP7_75t_R FILLER_46_24 ();
 DECAPx10_ASAP7_75t_R FILLER_46_46 ();
 DECAPx10_ASAP7_75t_R FILLER_46_68 ();
 DECAPx10_ASAP7_75t_R FILLER_46_90 ();
 DECAPx10_ASAP7_75t_R FILLER_46_112 ();
 DECAPx10_ASAP7_75t_R FILLER_46_134 ();
 DECAPx10_ASAP7_75t_R FILLER_46_156 ();
 DECAPx10_ASAP7_75t_R FILLER_46_178 ();
 DECAPx10_ASAP7_75t_R FILLER_46_200 ();
 DECAPx10_ASAP7_75t_R FILLER_46_222 ();
 DECAPx6_ASAP7_75t_R FILLER_46_244 ();
 DECAPx10_ASAP7_75t_R FILLER_47_2 ();
 DECAPx10_ASAP7_75t_R FILLER_47_24 ();
 DECAPx10_ASAP7_75t_R FILLER_47_46 ();
 DECAPx10_ASAP7_75t_R FILLER_47_68 ();
 DECAPx10_ASAP7_75t_R FILLER_47_90 ();
 DECAPx10_ASAP7_75t_R FILLER_47_112 ();
 DECAPx10_ASAP7_75t_R FILLER_47_134 ();
 DECAPx10_ASAP7_75t_R FILLER_47_156 ();
 DECAPx10_ASAP7_75t_R FILLER_47_178 ();
 DECAPx10_ASAP7_75t_R FILLER_47_200 ();
 DECAPx10_ASAP7_75t_R FILLER_47_222 ();
 DECAPx6_ASAP7_75t_R FILLER_47_244 ();
 DECAPx10_ASAP7_75t_R FILLER_48_2 ();
 DECAPx10_ASAP7_75t_R FILLER_48_24 ();
 DECAPx10_ASAP7_75t_R FILLER_48_46 ();
 DECAPx10_ASAP7_75t_R FILLER_48_68 ();
 DECAPx10_ASAP7_75t_R FILLER_48_90 ();
 DECAPx10_ASAP7_75t_R FILLER_48_112 ();
 DECAPx10_ASAP7_75t_R FILLER_48_134 ();
 DECAPx10_ASAP7_75t_R FILLER_48_156 ();
 DECAPx10_ASAP7_75t_R FILLER_48_178 ();
 DECAPx10_ASAP7_75t_R FILLER_48_200 ();
 DECAPx10_ASAP7_75t_R FILLER_48_222 ();
 DECAPx6_ASAP7_75t_R FILLER_48_244 ();
 DECAPx10_ASAP7_75t_R FILLER_49_2 ();
 DECAPx10_ASAP7_75t_R FILLER_49_24 ();
 DECAPx10_ASAP7_75t_R FILLER_49_46 ();
 DECAPx10_ASAP7_75t_R FILLER_49_68 ();
 DECAPx10_ASAP7_75t_R FILLER_49_90 ();
 DECAPx10_ASAP7_75t_R FILLER_49_112 ();
 DECAPx10_ASAP7_75t_R FILLER_49_134 ();
 DECAPx10_ASAP7_75t_R FILLER_49_156 ();
 DECAPx10_ASAP7_75t_R FILLER_49_178 ();
 DECAPx10_ASAP7_75t_R FILLER_49_200 ();
 DECAPx10_ASAP7_75t_R FILLER_49_222 ();
 DECAPx6_ASAP7_75t_R FILLER_49_244 ();
 DECAPx10_ASAP7_75t_R FILLER_50_2 ();
 DECAPx10_ASAP7_75t_R FILLER_50_24 ();
 DECAPx10_ASAP7_75t_R FILLER_50_46 ();
 DECAPx10_ASAP7_75t_R FILLER_50_68 ();
 DECAPx10_ASAP7_75t_R FILLER_50_90 ();
 DECAPx4_ASAP7_75t_R FILLER_50_112 ();
 FILLER_ASAP7_75t_R FILLER_50_122 ();
 DECAPx6_ASAP7_75t_R FILLER_50_129 ();
 DECAPx1_ASAP7_75t_R FILLER_50_143 ();
 DECAPx6_ASAP7_75t_R FILLER_50_152 ();
 DECAPx10_ASAP7_75t_R FILLER_50_176 ();
 DECAPx10_ASAP7_75t_R FILLER_50_198 ();
 DECAPx10_ASAP7_75t_R FILLER_50_220 ();
 DECAPx6_ASAP7_75t_R FILLER_50_242 ();
 FILLER_ASAP7_75t_R FILLER_50_256 ();
 DECAPx10_ASAP7_75t_R FILLER_51_2 ();
 DECAPx10_ASAP7_75t_R FILLER_51_24 ();
 DECAPx10_ASAP7_75t_R FILLER_51_46 ();
 DECAPx6_ASAP7_75t_R FILLER_51_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_82 ();
 DECAPx1_ASAP7_75t_R FILLER_51_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_102 ();
 DECAPx2_ASAP7_75t_R FILLER_51_108 ();
 FILLER_ASAP7_75t_R FILLER_51_114 ();
 DECAPx1_ASAP7_75t_R FILLER_51_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_125 ();
 DECAPx2_ASAP7_75t_R FILLER_51_136 ();
 FILLER_ASAP7_75t_R FILLER_51_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_144 ();
 DECAPx1_ASAP7_75t_R FILLER_51_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_159 ();
 FILLER_ASAP7_75t_R FILLER_51_165 ();
 DECAPx4_ASAP7_75t_R FILLER_51_177 ();
 DECAPx10_ASAP7_75t_R FILLER_51_192 ();
 DECAPx10_ASAP7_75t_R FILLER_51_214 ();
 DECAPx10_ASAP7_75t_R FILLER_51_236 ();
endmodule
